/*
Copyright (c) 2025 Kerim TURAK

Permission is granted to use, copy, modify, and distribute this software for any purpose,
with or without fee, provided that the above notice appears in all copies.

THE SOFTWARE IS PROVIDED "AS IS" WITHOUT ANY WARRANTY OF ANY KIND.
*/
`timescale 1ns / 1ps
`include "ceres_defines.svh"
module execution
  import ceres_param::*;
(
`ifdef COMMIT_TRACER
    output logic        [XLEN-1:0] csr_wr_data_o,
    output logic                   csr_write_valid_o,       // CSR write was accepted
`endif
    input  logic                   clk_i,
    input  logic                   rst_ni,
    input  stall_e                 stall_i,
    input  logic        [     1:0] fwd_a_i,
    input  logic        [     1:0] fwd_b_i,
    input  logic        [XLEN-1:0] alu_result_i,
    input  logic        [XLEN-1:0] wb_data_i,
    input  logic        [XLEN-1:0] r1_data_i,
    input  logic        [XLEN-1:0] r2_data_i,
    input  logic        [     1:0] alu_in1_sel_i,
    input  logic                   alu_in2_sel_i,
    input  logic                   rd_csr_i,
    input  logic                   wr_csr_i,
    input  logic        [    11:0] csr_idx_i,
    input  logic                   csr_or_data_i,
    input  logic                   trap_active_i,
    input  logic                   de_trap_active_i,
    input  logic        [XLEN-1:0] trap_cause_i,
    input  logic        [XLEN-1:0] trap_tval_i,             // faulting instruction / adres
    input  logic        [XLEN-1:0] trap_mepc_i,
    // Hardware interrupt inputs
    input  logic                   timer_irq_i,             // CLINT timer interrupt
    input  logic                   sw_irq_i,                // CLINT software interrupt
    input  logic                   ext_irq_i,               // PLIC external interrupt
    input  logic        [XLEN-1:0] pc_i,
    input  logic        [XLEN-1:0] pc_incr_i,
    input  logic        [XLEN-1:0] imm_i,
    input  pc_sel_e                pc_sel_i,
    input  alu_op_e                alu_ctrl_i,
    input  instr_type_e            instr_type_i,
    input  logic                   misa_c_i,                // C extension state when instruction was fetched
    output logic        [XLEN-1:0] write_data_o,
    output logic        [XLEN-1:0] pc_target_o,
    output logic        [XLEN-1:0] alu_result_o,
    output logic                   pc_sel_o,
    output logic                   alu_stall_o,
    output exc_type_e              exc_type_o,
    output logic        [XLEN-1:0] mtvec_o,
    output logic                   misa_c_o,
    output logic        [XLEN-1:0] tdata1_o         [0:1],
    output logic        [XLEN-1:0] tdata2_o         [0:1],
    output logic        [XLEN-1:0] tcontrol_o

);

  logic        [XLEN-1:0] data_a;
  logic        [XLEN-1:0] operant_a;
  logic        [XLEN-1:0] operant_b;
  logic signed [XLEN-1:0] signed_imm;
  logic                   ex_zero;
  logic                   ex_slt;
  logic                   ex_sltu;
  logic        [XLEN-1:0] tdata1             [0:1];
  logic        [XLEN-1:0] tdata2             [0:1];
  logic        [XLEN-1:0] tcontrol;
  logic        [XLEN-1:0] alu_result;
  logic        [XLEN-1:0] csr_rdata;
  logic        [XLEN-1:0] mepc;
  logic                   misa_c;
  logic        [XLEN-1:0] tcontrol_effective;
  logic        [XLEN-1:0] tdata1_effective   [0:1];
  logic        [XLEN-1:0] tdata2_effective   [0:1];
  logic                   trigger0_hit;
  logic                   trigger1_hit;
  logic                   target_misaligned;
  assign misa_c_o = misa_c;

  always_comb begin
    data_a = fwd_a_i[1] ? alu_result_i : (fwd_a_i[0] ? wb_data_i : r1_data_i);
    case (alu_in1_sel_i)
      2'b00: operant_a = data_a;
      2'b01: operant_a = pc_incr_i;
      2'b10: operant_a = pc_i;
      2'b11: operant_a = data_a;
    endcase

    write_data_o = fwd_b_i[1] ? alu_result_i : (fwd_b_i[0] ? wb_data_i : r2_data_i);
    operant_b = alu_in2_sel_i ? imm_i : write_data_o;
    signed_imm = imm_i;
    /*
    Eğer exception desteği yoksa burası
    pc_target_o = pc_sel_i == JALR ? (data_a + imm_i) & ~1 : pc_i + signed_imm;
    */
    pc_target_o = instr_type_i == mret ? mepc : pc_sel_i == JALR ? (data_a + imm_i) & ~1 : pc_i + signed_imm;

    pc_sel_o = (pc_sel_i == BEQ) && ex_zero;
    pc_sel_o |= (pc_sel_i == BNE) && !ex_zero;
    pc_sel_o |= (pc_sel_i == BLT) && ex_slt;
    pc_sel_o |= (pc_sel_i == BGE) && (!ex_slt || ex_zero);
    pc_sel_o |= (pc_sel_i == BLTU) && ex_sltu;
    pc_sel_o |= (pc_sel_i == BGEU) && (!ex_sltu || ex_zero);
    pc_sel_o |= (pc_sel_i == JALR);
    pc_sel_o |= (pc_sel_i == JAL);
    pc_sel_o |= (instr_type_i == mret);

    // ------------------------------------------------------------------------
    // LOCAL CSR WRITE BYPASS for same-cycle breakpoint detection
    // ------------------------------------------------------------------------
    // When writing to trigger CSRs, use alu_result directly to enable
    // immediate breakpoint detection without waiting for next cycle.
    // This local bypass does NOT create combinational loop because:
    // - It's local to execution stage (doesn't feedback through trap_active)
    // - CSR file outputs are registered (tcontrol_out_reg breaks the loop)


    tcontrol_effective = (wr_csr_i && csr_idx_i == 12'h7A5) ? alu_result : tcontrol;
    // Trigger 0 bypass
    tdata1_effective[0] = (wr_csr_i && csr_idx_i == 12'h7A1) ? alu_result : tdata1[0];
    tdata2_effective[0] = (wr_csr_i && csr_idx_i == 12'h7A2) ? alu_result : tdata2[0];
    // Trigger 1 bypass
    tdata1_effective[1] = (wr_csr_i && csr_idx_i == 12'h7A1) ? alu_result : tdata1[1];
    tdata2_effective[1] = (wr_csr_i && csr_idx_i == 12'h7A2) ? alu_result : tdata2[1];

    // LOAD/STORE breakpoint detection for both triggers
    // tdata1[0] = LOAD match enable, tdata1[1] = STORE match enable
    // tdata1[6] = M-mode match, tdata1[31:28] = type (2 = mcontrol)
    // tcontrol[3] = MTE (M-mode Trigger Enable)

    // Check Trigger 0
    trigger0_hit = 1'b0;
    if (tcontrol_effective[3] && tdata1_effective[0][6] && (tdata1_effective[0][31:28] == 4'h2)) begin
      if (tdata1_effective[0][0] && (instr_type_i inside {i_lb, i_lh, i_lw, i_lbu, i_lhu})) begin
        trigger0_hit = (alu_result == tdata2_effective[0]);
      end else if (tdata1_effective[0][1] && (instr_type_i inside {s_sb, s_sh, s_sw})) begin
        trigger0_hit = (alu_result == tdata2_effective[0]);
      end
    end

    // Check Trigger 1
    trigger1_hit = 1'b0;
    if (tcontrol_effective[3] && tdata1_effective[1][6] && (tdata1_effective[1][31:28] == 4'h2)) begin
      if (tdata1_effective[1][0] && (instr_type_i inside {i_lb, i_lh, i_lw, i_lbu, i_lhu})) begin
        trigger1_hit = (alu_result == tdata2_effective[1]);
      end else if (tdata1_effective[1][1] && (instr_type_i inside {s_sb, s_sh, s_sw})) begin
        trigger1_hit = (alu_result == tdata2_effective[1]);
      end
    end

    // Jump/Branch target misalignment check:
    // - If C extension enabled (misa_c=1): target must be 2-byte aligned (pc_target[0]=0)
    // - If C extension disabled (misa_c=0): target must be 4-byte aligned (pc_target[1:0]=00)
    // IMPORTANT: Use misa_c_i (pipelined value from when instruction was fetched)
    // instead of misa_c (current CSR value) to handle MISA.C changes in flight
    if (misa_c_i) begin
      target_misaligned = pc_target_o[0];  // 2-byte alignment check
    end else begin
      target_misaligned = (pc_target_o[1:0] != 2'b00);  // 4-byte alignment check
    end

    // Priority: Trigger hit > Instruction misaligned
    // Exception check priority:
    // 1. Hardware breakpoint (trigger)
    // 2. Jump/Branch target misalignment
    // Note: MRET target (mepc) is exempt from alignment check because mepc is
    // aligned when written. This prevents spurious exceptions when MISA.C changes
    // between trap entry and return.
    if (trigger0_hit || trigger1_hit) begin
      exc_type_o = BREAKPOINT;
    end else if (instr_type_i == mret) begin
      exc_type_o = NO_EXCEPTION;  // MRET: mepc already aligned when written
    end else begin
      exc_type_o = pc_sel_o && target_misaligned ? INSTR_MISALIGNED : NO_EXCEPTION;
    end
  end

  alu i_alu (
      .clk_i      (clk_i),
      .rst_ni     (rst_ni),
      .alu_a_i    (operant_a),
      .csr_rdata_i(csr_rdata),
      .alu_b_i    (operant_b),
      .op_sel_i   (alu_ctrl_i),
      .alu_stall_o(alu_stall_o),
      .zero_o     (ex_zero),
      .slt_o      (ex_slt),
      .sltu_o     (ex_sltu),
      .alu_o      (alu_result)
  );

  logic [XLEN-1:0] rd_data;

  always_comb begin
    unique case (instr_type_i)
      u_jal, i_jalr: rd_data = pc_incr_i;  // rd = PC+4
      default:       rd_data = alu_result;
    endcase

    if (rd_csr_i && csr_or_data_i) rd_data = csr_rdata;
  end

  assign alu_result_o = rd_data;

`ifdef COMMIT_TRACER
  always_comb begin
    if (instr_type_i == mret) begin
      // cs_reg_file içindeki pack_mstatus sonucu loglanmalı
      csr_wr_data_o        = 0;
      csr_wr_data_o[3]     = csr_rdata[3];
      csr_wr_data_o[7]     = csr_rdata[7];
      csr_wr_data_o[12:11] = csr_rdata[12:11];
    end else begin
      csr_wr_data_o = csr_wmask(csr_idx_i, alu_result);
    end
  end
`endif

  cs_reg_file i_cs_reg_file (
      .clk_i            (clk_i),
      .rst_ni           (rst_ni),
      .stall_i          (stall_i),
      .rd_en_i          (rd_csr_i),
      .wr_en_i          (wr_csr_i),
      .csr_idx_i        (csr_idx_i),
      .csr_wdata_i      (alu_result),
      .csr_rdata_o      (csr_rdata),
      .trap_active_i    (trap_active_i),
      .de_trap_active_i (de_trap_active_i),
      .trap_cause_i     (trap_cause_i),
      .trap_mepc_i      (trap_mepc_i),
      .trap_tval_i      (trap_tval_i),
      .pc_i             (pc_i),
      .instr_type_i     (instr_type_i),
      // Hardware interrupt inputs
      .timer_irq_i      (timer_irq_i),
      .sw_irq_i         (sw_irq_i),
      .ext_irq_i        (ext_irq_i),
      .mtvec_o          (mtvec_o),
      .mepc_o           (mepc),
      .misa_c_o         (misa_c),
`ifdef COMMIT_TRACER
      .csr_write_valid_o(csr_write_valid_o),
`endif
      .tdata1_o         (tdata1),
      .tdata2_o         (tdata2),
      .tcontrol_o       (tcontrol)
  );

  assign tdata1_o   = tdata1;
  assign tdata2_o   = tdata2;
  assign tcontrol_o = tcontrol;
endmodule
