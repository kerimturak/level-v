@80000000
97 31 00 00 93 81 C1 1F 17 01 01 00 13 01 81 FF
97 32 00 00 93 82 02 1F 17 33 00 00 13 03 43 20
63 86 62 00 23 A0 02 00 91 02 DD BF 93 02 00 00
63 83 02 00 82 92 97 02 00 00 93 82 22 6B 63 83
02 00 82 92 01 A0
@80000046
19 C6 03 15 25 00 83 97 25 00 1D 8D 82 80 83 17
05 00 93 96 07 01 13 F7 07 F0 93 D7 86 01 D9 8F
23 10 F5 00 83 97 05 00 03 15 25 00 93 96 07 01
13 F7 07 F0 93 D7 86 01 D9 8F 23 90 F5 00 83 97
25 00 1D 8D 82 80 03 18 05 00 93 57 78 40 85 8B
81 C7 13 75 F8 07 82 80 13 57 38 40 3D 8B 01 11
93 17 47 00 33 06 F7 00 22 CC 06 CE 26 CA 93 76
78 00 83 D7 85 03 AE 88 2A 84 32 87 B5 C6 05 46
63 9F C6 04 3E 86 13 85 88 02 BA 85 42 C6 46 C4
EF 10 20 0C A2 48 93 14 05 01 32 48 83 D7 C8 03
C1 84 BD EF 83 D7 88 03 23 9E A8 02 BE 85 46 C6
42 C4 EF 10 E0 5D 22 48 B2 48 AA 87 13 78 08 F0
13 F5 F4 07 33 68 05 01 23 9C F8 02 13 68 08 08
F2 40 23 10 04 01 62 44 D2 44 05 61 82 80 13 15
08 01 41 81 C2 84 D9 B7 93 06 10 02 63 E4 C6 00
13 07 20 02 83 96 28 00 03 96 08 00 83 A5 48 01
03 A5 88 01 42 C6 46 C4 EF 10 C0 34 A2 48 93 14
05 01 32 48 83 D7 E8 03 C1 84 99 E3 23 9F A8 02
83 D7 88 03 61 B7 01 11 26 CA AE 84 B2 85 06 CE
22 CC 32 C6 09 3F B2 45 2A 84 26 85 29 37 F2 40
33 05 A4 40 62 44 D2 44 05 61 82 80 03 97 05 00
83 97 25 00 23 10 E5 00 23 11 F5 00 82 80 03 28
06 00 93 08 88 00 63 FF E8 02 98 42 13 03 47 00
63 7A F3 02 23 20 16 01 1C 41 83 98 05 00 03 96
25 00 23 20 F8 00 23 20 05 01 23 22 E8 00 9C 42
42 85 91 07 9C C2 83 27 48 00 23 90 17 01 23 91
C7 00 82 80 01 48 42 85 82 80 AA 87 08 41 D4 43
50 41 18 41 D0 C3 54 C1 98 C3 23 20 05 00 82 80
D4 41 58 41 9C 41 54 C1 D8 C1 1C C1 88 C1 82 80
03 97 25 00 63 4C 07 00 01 E5 82 80 08 41 15 C1
5C 41 83 97 27 00 E3 9B E7 FE 82 80 19 C9 03 97
05 00 19 A0 08 41 11 C5 5C 41 83 C7 07 00 E3 9B
E7 FE 82 80 01 C9 01 47 11 A0 3E 85 1C 41 18 C1
2A 87 E5 FF 82 80 79 71 4A D0 56 CA 5A C8 5E C6
6A C0 85 4A 06 D6 22 D4 26 D2 4E CE 52 CC 62 C4
66 C2 2A 89 AE 8B 32 8B 56 8D 63 01 09 0A 81 4C
81 44 01 4C 85 0C CA 87 01 44 63 55 54 01 9C 43
05 04 E5 FF CA 89 56 8A 3E 89 63 5F 80 00 63 04
0A 00 63 11 09 02 A6 87 7D 14 CE 84 83 A9 09 00
85 CB 84 C3 E3 45 80 FE B3 37 20 01 63 57 40 05
B1 C7 05 C8 83 25 49 00 03 A5 49 00 5A 86 82 9B
63 59 A0 04 A6 87 7D 1A CA 84 03 29 09 00 F1 FB
26 8C 65 BF 98 C0 B3 37 20 01 BA 84 63 0E 0A 00
81 CF 4A 87 7D 1A 03 29 09 00 ED F4 3A 8C B3 37
20 01 BA 84 E3 16 0A FE BA 84 AD FF 23 A0 04 00
63 88 AC 03 62 89 86 0A E3 13 09 F6 23 20 00 00
02 90 03 A7 09 00 7D 14 91 C4 A6 87 CE 84 84 C3
BA 89 49 B7 4E 8C CE 84 BA 89 E3 45 80 F8 AD BF
B2 50 22 54 92 54 02 59 F2 49 62 4A D2 4A 42 4B
B2 4B 92 4C 02 4D 62 85 22 4C 45 61 82 80 03 16
45 00 79 71 22 D4 06 D6 26 D2 4A D0 4E CE 40 51
63 5D C0 1C 63 CF 05 1C 63 06 04 1E AE 86 01 4E
01 4F 81 4E 81 48 01 43 A2 87 19 A0 9C 43 C9 CF
D8 43 03 18 27 00 E3 1B D8 FE 81 46 11 A0 3A 84
18 40 14 C0 A2 86 65 FF D1 C3 D8 43 85 0E 03 17
07 00 93 76 17 00 81 C6 25 87 05 8B BA 98 98 43
11 C7 14 43 94 C3 1C 40 1C C3 18 C0 63 48 08 02
93 07 1E 00 13 9E 07 01 93 06 18 00 C2 06 C2 07
13 5E 0E 41 C1 86 C1 83 63 0D C6 05 13 F3 F7 0F
E3 DC 06 F8 9A 86 A2 87 61 78 0D A0 93 06 1E 00
13 9E 06 01 13 5E 0E 41 C2 06 C1 82 63 0A C6 03
93 F6 F6 0F A2 87 19 A0 9C 43 8D C3 D8 43 03 43
07 00 E3 1B D3 FE 95 BF 36 88 85 BF 1C 40 05 0F
DC 43 83 87 17 00 85 8B BE 98 49 BF 36 83 B1 BF
C2 86 93 97 2E 00 B3 87 E7 41 BE 98 93 94 08 01
C1 80 63 5E B0 00 2A 86 97 05 00 00 93 85 E5 D0
22 85 1A C6 36 C4 C5 3B 32 43 A2 46 2A 84 1C 40
22 89 83 A9 07 00 D8 43 83 A5 49 00 03 A6 09 00
CC C3 23 A2 E9 00 90 C3 23 A0 09 00 63 D7 06 00
71 A0 03 29 09 00 63 0A 09 08 83 27 49 00 83 97
27 00 E3 98 D7 FE 5C 40 A6 85 03 95 07 00 EF 10
00 72 03 29 09 00 AA 84 E3 17 09 FE 03 29 04 00
03 A7 49 00 83 26 49 00 83 27 09 00 22 85 23 A2
D9 00 23 22 E9 00 23 A0 F9 00 23 20 39 01 01 46
97 05 00 00 93 85 05 B6 BD 33 00 41 2A 89 19 C8
83 27 49 00 A6 85 03 95 07 00 EF 10 40 6D 00 40
AA 84 7D F4 B2 50 22 54 02 59 F2 49 26 85 92 54
45 61 82 80 03 29 09 00 63 09 09 00 83 27 49 00
83 C7 07 00 E3 18 F3 FE BD BF 03 29 04 00 E3 0B
09 F8 5C 40 A6 85 03 95 07 00 EF 10 40 69 03 29
09 00 AA 84 E3 11 09 F6 95 BF AE 86 81 44 01 43
09 B7 09 C8 2E 88 A2 87 81 48 81 46 01 4F 01 4E
81 4E 6D BD 81 47 9C 43 02 90 B7 D7 CC CC 93 87
D7 CC 33 35 F5 02 E1 77 23 A0 05 00 93 87 07 08
93 86 05 01 13 83 85 00 61 77 11 81 93 08 E5 FF
13 9E 38 00 2E 9E 23 A2 C5 01 23 10 FE 00 13 9F
28 00 23 11 0E 00 72 9F 93 07 4E 00 63 FA C6 0D
13 08 8E 00 63 76 E8 0D DC C5 23 A4 05 00 23 A0
65 00 13 47 F7 FF FD 57 23 13 EE 00 23 12 FE 00
E1 7F 93 CF FF FF 01 47 63 85 08 04 B3 47 C7 00
8E 07 13 75 77 00 93 F7 87 07 C9 8F 93 9E 87 00
13 83 86 00 05 07 13 05 48 00 F6 97 63 71 C3 03
63 7F E5 01 83 AE 05 00 23 A0 D6 01 94 C1 23 A2
06 01 23 10 F8 00 23 11 F8 01 9A 86 2A 88 E3 9F
E8 FA 88 41 14 41 B1 C6 B7 D7 CC CC 93 87 D7 CC
B3 B8 F8 02 11 6E 7D 1E 13 08 00 20 05 47 93 D8
28 00 11 A0 9A 86 93 77 08 70 33 43 E6 00 B3 E7
67 00 48 41 B3 F7 C7 01 63 73 17 01 BA 87 03 A3
06 00 23 11 F5 00 05 07 13 08 08 10 36 85 E3 1B
03 FC 2E 85 01 46 97 05 00 00 93 85 A5 9C E1 BE
3E 88 9A 86 B1 B7 41 11 4A C0 03 29 C5 01 06 C6
23 2C 05 02 23 2E 05 02 63 00 09 04 22 C4 26 C2
2A 84 81 44 85 45 22 85 5D 39 83 55 84 03 EF 10
20 02 23 1C A4 02 FD 55 22 85 55 31 83 55 84 03
EF 10 00 01 23 1C A4 02 99 E0 23 1D A4 02 85 04
E3 1A 99 FC 22 44 92 44 B2 40 02 49 01 45 41 01
82 80 59 71 86 D6 A2 D4 A6 D2 CA D0 CE CE D2 CC
D6 CA DA C8 DE C6 E2 C4 E6 C2 EA C0 13 01 01 81
2E 86 2A C6 6C 00 13 05 E1 05 EF 10 20 71 05 45
EF 00 50 69 23 1E A1 00 09 45 EF 00 B0 68 23 1F
A1 00 0D 45 EF 00 10 68 23 10 A1 02 11 45 EF 00
70 67 2A DC 15 45 13 04 01 83 EF 00 B0 66 11 E1
1D 45 2A DE 83 27 C4 7E 63 8F 07 24 05 47 63 8F
E7 4E 93 77 25 00 B3 37 F0 00 13 03 01 06 13 77
15 00 3E 97 23 1E 01 04 23 2A 64 7E 93 77 45 00
81 C7 05 07 42 07 41 83 93 05 00 7D B3 D5 E5 02
64 08 A6 86 81 47 01 46 85 48 0D 48 2E DA 33 97
F8 00 69 8F 85 07 63 1E 07 0E 91 06 E3 99 07 FF
F2 57 13 F7 17 00 09 CB 03 16 C4 7E 83 25 84 7F
52 55 65 3B F2 57 AA C0 13 F7 27 00 55 EF 91 8B
99 C7 42 56 83 15 C4 7E 52 55 EF 00 90 1E E2 57
85 EF 85 47 3E DC 62 57 93 17 27 00 BA 97 86 07
3E DC EF 10 80 5B 26 85 79 3D EF 10 60 5D EF 10
80 5F EF 10 A0 61 65 D1 A9 47 B3 D7 A7 02 62 57
85 07 B3 87 E7 02 3E DC EF 10 20 59 26 85 A5 3D
EF 10 00 5B EF 10 20 5D AA 89 03 15 C4 7E AE 8A
81 45 EF 10 C0 3A AA 85 03 15 E4 7E EF 10 20 3A
AA 85 03 15 04 7F EF 10 80 39 AA 85 03 15 41 03
EF 10 E0 38 A1 67 93 87 57 B0 2A 8A 63 00 F5 3E
63 F9 A7 04 A5 67 93 87 27 A0 63 01 F5 3C BD 67
93 87 57 9F 63 1A F5 14 17 25 00 00 13 05 A5 FD
EF 10 10 06 8D 47 B9 A0 83 17 E4 7E 03 16 C4 7E
83 25 C4 7F 52 55 C2 07 5D 8E D4 00 ED 26 F2 57
3D B7 33 07 B6 02 05 06 42 06 41 82 1A 97 D8 C6
ED BD 89 67 93 87 27 8F 63 0A F5 38 95 67 93 87
F7 EA 63 13 F5 10 17 25 00 00 13 05 85 F5 EF 10
30 01 89 47 97 3B 00 00 93 8B 6B 92 03 A7 0B 00
63 0D 07 38 86 07 17 2D 00 00 13 0D 8D 48 3E 9D
81 4C 01 4B 05 6C 1D A0 B3 87 64 01 8A 07 A2 97
E2 97 83 D7 C7 82 33 89 97 01 05 0B 83 A7 0B 00
42 0B 13 5B 0B 01 CA 8C 63 7F FB 0A 93 14 4B 00
33 89 64 01 0A 09 22 99 62 99 83 27 C9 80 23 16
09 82 13 F7 17 00 0D C7 03 56 69 82 83 56 0D 00
63 00 D6 02 DA 85 17 25 00 00 13 05 85 F6 EF 10
20 79 03 57 C9 82 83 27 C9 80 05 07 23 16 E9 82
13 F7 27 00 15 CB 33 89 64 01 0A 09 22 99 62 99
03 56 89 82 83 56 CD 00 63 00 D6 02 DA 85 17 25
00 00 13 05 05 F6 EF 10 A0 75 03 57 C9 82 83 27
C9 80 05 07 23 16 E9 82 91 8B B9 DF DA 94 8A 04
A2 94 E2 94 03 D6 A4 82 83 56 8D 01 63 18 D6 20
83 D7 C4 82 89 BF 83 17 04 7F E3 94 07 DA 93 07
60 06 23 18 F4 7E 71 BB C1 67 13 89 F7 FF 97 3B
00 00 93 8B CB 82 EF 10 C0 3A D2 55 2A 99 17 25
00 00 13 05 45 F6 EF 10 A0 6F CE 85 17 25 00 00
13 05 E5 F6 EF 10 C0 6E D6 85 4E 85 EF 10 00 42
AA 85 17 25 00 00 13 05 05 F7 EF 10 60 6D 4E 85
D6 85 EF 10 A0 40 63 1A 05 1C 4E 85 D6 85 EF 10
E0 3F A5 47 63 FB A7 1A 83 A7 0B 00 E2 55 17 25
00 00 13 05 45 FB 42 09 B3 85 F5 02 13 59 09 41
EF 10 00 6A 97 25 00 00 93 85 65 FB 17 25 00 00
13 05 A5 FB EF 10 C0 68 97 25 00 00 93 85 65 FC
17 25 00 00 13 05 65 06 EF 10 80 67 97 25 00 00
93 85 25 07 17 25 00 00 13 05 25 07 EF 10 40 66
D2 85 17 25 00 00 13 05 C5 07 EF 10 60 65 F2 57
13 F7 17 00 0D CF 03 A7 0B 00 15 CB 81 44 85 69
93 97 44 00 A6 97 8A 07 A2 97 CE 97 03 D6 67 82
A6 85 17 25 00 00 13 05 85 06 EF 10 60 62 85 04
83 A7 0B 00 C2 04 C1 80 E3 EC F4 FC F2 57 13 F7
27 00 15 CF 03 A7 0B 00 63 03 07 1A 81 44 85 69
93 97 44 00 A6 97 8A 07 A2 97 CE 97 03 D6 87 82
A6 85 17 25 00 00 13 05 45 04 EF 10 60 5E 85 04
83 A7 0B 00 C2 04 C1 80 E3 EC F4 FC F2 57 91 8B
85 CF 83 A7 0B 00 81 44 85 69 B5 C3 93 97 44 00
A6 97 8A 07 A2 97 CE 97 03 D6 A7 82 A6 85 17 25
00 00 13 05 45 02 EF 10 A0 5A 85 04 83 A7 0B 00
C2 04 C1 80 E3 EC F4 FC 83 A7 0B 00 81 44 85 69
9D C7 93 97 44 00 A6 97 8A 07 A2 97 CE 97 03 D6
47 82 A6 85 17 25 00 00 13 05 A5 00 EF 10 40 57
85 04 83 A7 0B 00 C2 04 C1 80 E3 EC F4 FC 63 09
09 08 63 5E 20 09 17 25 00 00 13 05 45 0B EF 10
20 55 13 05 E1 05 EF 10 A0 2A 13 01 01 7F B6 50
26 54 96 54 06 59 F6 49 66 4A D6 4A 46 4B B6 4B
26 4C 96 4C 06 4D 01 45 65 61 82 80 DA 85 17 25
00 00 13 05 45 D5 EF 10 A0 51 83 D7 C4 82 85 07
C2 07 C1 83 23 96 F4 82 3D B3 17 25 00 00 13 05
85 DC EF 10 E0 4F 05 09 81 B5 E2 54 83 A7 0B 00
D6 85 4E 85 B3 84 F4 02 EF 10 40 22 AA 85 17 25
00 00 13 05 C5 D8 B3 D5 B4 02 EF 10 60 4D 31 B5
17 25 00 00 13 05 A5 F7 EF 10 80 4C 9D BF 17 25
00 00 13 05 85 FB EF 10 A0 4B A5 B7 17 25 00 00
13 05 65 B9 EF 10 C0 4A 81 47 69 B9 17 25 00 00
13 05 65 BB EF 10 C0 49 85 47 69 B1 17 25 00 00
13 05 65 C3 EF 10 C0 48 91 47 AD B9 83 17 04 7F
E3 91 07 B0 B7 37 15 34 93 87 57 41 13 07 60 06
23 26 F4 7E 23 18 E4 7E ED B4 01 49 A9 BB 91 8B
E3 84 07 EC ED BD 41 11 22 C6 26 C4 2A 88 11 E2
05 46 13 84 F5 FF 71 98 93 03 44 00 81 47 63 0B
08 08 3E 85 85 07 33 87 F7 02 0E 07 E3 6B 07 FF
B3 02 A5 02 86 02 33 84 53 00 59 C1 4A C2 AA 84
13 03 15 00 13 19 15 00 22 8F 81 4E 85 47 33 8E
83 40 BE 8F FA 85 33 06 F6 02 B3 08 BE 00 89 05
13 57 F6 41 41 83 3A 96 42 06 41 82 19 8E 33 88
C7 00 33 07 F8 00 23 9F 05 FF 13 77 F7 0F 85 07
23 90 E8 00 E3 99 67 FC 85 0E B3 07 F5 01 2A 93
4A 9F E3 90 AE FC 12 49 B3 07 54 00 FD 17 80 C6
F1 9B 32 44 91 07 84 C2 DC C6 23 A2 76 00 A2 44
41 01 82 80 FD 54 4A C2 19 04 26 85 89 42 49 B7
81 42 81 44 D1 BF AA 8E 29 C9 13 1E 25 00 B3 88
C5 01 01 43 01 45 01 47 81 46 B3 87 C8 41 09 A8
33 08 B5 00 13 15 08 01 91 07 41 85 63 82 F8 02
BA 85 98 43 13 08 A5 00 BA 96 B3 A5 E5 00 E3 51
D6 FE 13 15 08 01 91 07 81 46 41 85 E3 92 F8 FE
05 03 F2 98 E3 93 6E FC 82 80 01 45 82 80 1D C9
13 1E 15 00 33 08 C6 01 01 43 81 48 13 16 23 00
2E 96 B3 07 C8 41 03 97 07 00 89 07 11 06 33 07
D7 02 23 2E E6 FE E3 18 F8 FE 85 08 2A 93 72 98
E3 1E 15 FD 82 80 05 C5 13 18 15 00 B3 86 05 01
81 45 B3 87 06 41 03 D7 07 00 89 07 32 97 23 9F
E7 FE E3 9A F6 FE 85 05 C2 96 E3 14 B5 FE 82 80
15 CD 13 1F 25 00 13 1E 15 00 2E 9F 36 9E 81 4E
13 98 1E 00 32 98 B6 87 81 48 03 17 08 00 03 93
07 00 89 07 09 08 33 07 67 02 BA 98 E3 17 FE FE
23 A0 15 01 91 05 AA 9E E3 1C BF FC 82 80 35 C1
41 11 13 13 15 00 22 C6 B2 82 36 84 33 0E 66 00
81 43 81 46 93 9E 23 00 AE 9E 22 8F 81 4F 7A 86
96 87 01 48 03 97 07 00 83 18 06 00 89 07 1A 96
33 07 17 03 3A 98 E3 17 FE FE 23 A0 0E 01 93 87
1F 00 91 0E 09 0F 63 04 F5 00 BE 8F C9 BF 9A 92
AA 93 1A 9E 63 84 F6 01 85 06 6D BF 32 44 41 01
82 80 82 80 35 C9 41 11 13 13 15 00 22 C6 B2 82
36 84 33 0E 66 00 81 43 81 46 93 9E 23 00 AE 9E
22 8F 81 4F 7A 88 16 86 81 48 03 17 08 00 83 17
06 00 09 06 1A 98 B3 87 E7 02 13 D7 27 40 95 87
3D 8B 93 F7 F7 07 B3 07 F7 02 BE 98 E3 1F CE FC
23 A0 1E 01 93 87 1F 00 91 0E 09 0F 63 04 F5 00
BE 8F C9 B7 9A 92 AA 93 1A 9E 63 84 F6 01 85 06
6D B7 32 44 41 01 82 80 82 80 79 71 4A D0 4E CE
56 CA 06 D6 22 D4 AE 8A 32 89 B6 89 63 09 05 22
93 15 15 00 26 D2 52 CC 2E 96 3A 8A FD 74 5A C8
5E C6 62 C4 66 C2 32 87 B3 64 9A 00 01 4B B3 07
B7 40 83 D6 07 00 89 07 D2 96 23 9F D7 FE E3 9A
E7 FE 13 04 1B 00 33 87 B7 00 63 04 85 00 22 8B
F9 BF 01 45 01 48 13 17 25 00 56 97 B3 07 B6 40
83 96 07 00 89 07 11 07 B3 86 46 03 23 2E D7 FE
E3 18 F6 FE 22 95 2E 96 63 04 68 01 05 08 E1 BF
13 1C 24 00 B3 8B 8A 01 5E 88 81 46 01 47 01 45
81 48 B3 07 88 41 09 A8 B3 05 C5 00 13 95 05 01
91 07 41 85 63 02 F8 02 36 86 94 43 93 05 A5 00
36 97 33 26 D6 00 E3 D1 E4 FE 13 95 05 01 91 07
01 47 41 85 E3 12 F8 FE 62 98 63 04 1B 01 85 08
C9 B7 81 45 EF 00 B0 3E CE 86 AA 8C 4A 86 22 85
D6 85 FD 3B 81 46 01 47 01 45 01 48 B3 87 8B 41
09 A8 B3 05 C5 00 13 95 05 01 91 07 41 85 63 82
77 03 36 86 94 43 93 05 A5 00 36 97 33 26 D6 00
E3 D1 E4 FE 13 95 05 01 91 07 01 47 41 85 E3 92
77 FF B3 8B 87 01 63 04 68 01 05 08 C1 B7 E6 85
EF 00 F0 38 CE 86 2A 8B 4A 86 22 85 D6 85 C5 33
01 43 81 47 81 46 01 45 81 48 13 16 23 00 56 96
81 45 11 A8 33 08 E5 00 13 15 08 01 85 05 41 85
11 06 63 F3 85 02 3E 87 1C 42 13 08 A5 00 BE 96
33 27 F7 00 E3 D0 D4 FE 13 15 08 01 85 05 81 46
41 85 11 06 E3 E1 85 FE 85 08 22 93 E3 EF 88 FA
DA 85 EF 00 D0 32 CE 86 2A 8B 4A 86 22 85 D6 85
D5 33 01 43 81 47 81 46 01 45 81 48 13 16 23 00
56 96 81 45 11 A8 33 08 E5 00 13 15 08 01 85 05
41 85 11 06 63 F3 85 02 3E 87 1C 42 13 08 A5 00
BE 96 33 27 F7 00 E3 D0 D4 FE 13 15 08 01 85 05
81 46 41 85 11 06 E3 E1 85 FE 85 08 22 93 E3 EF
88 FA DA 85 EF 00 B0 2C 81 45 01 46 93 97 15 00
CA 97 01 47 83 D6 07 00 05 07 89 07 B3 86 46 41
23 9F D7 FE E3 68 87 FE 05 06 A2 95 E3 60 86 FE
92 54 62 4A 42 4B B2 4B 22 4C 92 4C B2 50 22 54
42 05 02 59 F2 49 D2 4A 41 85 45 61 82 80 81 45
EF 00 F0 27 CE 86 4A 86 2A 84 D6 85 01 45 49 39
A2 85 01 45 EF 00 B0 26 CE 86 4A 86 2A 84 D6 85
01 45 75 39 A2 85 01 45 EF 00 70 25 2A 84 D6 85
CE 86 4A 86 01 45 39 33 A2 85 01 45 EF 00 30 24
75 B7 41 11 22 C4 14 45 32 84 2E 87 50 41 4C 45
08 41 06 C6 9D 33 A2 85 22 44 B2 40 41 01 6F 00
10 22 93 08 F5 FF 85 4E 63 F3 1E 0D F6 95 C2 05
C1 81 41 11 13 98 B5 01 22 C6 1D 43 93 F6 75 00
01 47 17 2E 00 00 13 0E 0E BB 11 4F 93 0F C0 02
93 57 E8 01 63 8E 66 04 63 66 DF 08 F5 16 C2 06
8A 07 C1 82 F2 97 63 EC DE 06 9C 4B A1 42 93 06
17 00 33 84 56 00 63 77 14 05 85 05 32 97 C2 05
C1 81 BA 86 B3 83 57 00 03 C8 07 00 85 07 85 06
A3 8F 06 FF E3 9A F3 FE 16 97 23 00 F7 01 13 98
B5 01 93 F6 75 00 22 87 93 57 E8 01 E3 96 66 FA
8A 07 A1 42 93 06 17 00 F2 97 33 84 56 00 9C 5B
E3 6D 14 FB 63 64 A7 00 01 A8 85 06 32 97 23 00
07 00 36 87 E3 EB A6 FE 32 44 41 01 82 80 9C 43
91 42 71 B7 8A 07 F2 97 9C 53 A1 42 49 B7 F6 86
01 47 11 A0 85 06 32 97 23 00 07 00 36 87 E3 EB
A6 FE 82 80 14 41 83 C7 06 00 8D CB 13 07 C0 02
63 8A E7 16 13 08 E0 02 63 8B 07 15 63 63 F8 02
93 87 57 FD 93 F7 D7 0F 63 81 07 16 D8 41 9C 41
85 06 05 07 85 07 9C C1 D8 C1 85 47 14 C1 3E 85
82 80 93 87 07 FD 93 F7 F7 0F 25 46 E3 60 F6 FE
90 41 93 87 16 00 05 06 90 C1 83 C6 16 00 63 82
06 16 63 87 E6 16 13 07 E0 02 63 8B E6 02 93 86
06 FD 93 F6 F6 0F 25 47 63 7C D7 00 98 49 93 86
17 00 85 47 3E 97 98 C9 14 C1 3E 85 82 80 90 C5
83 C6 17 00 85 07 63 86 06 12 13 07 C0 02 D1 B7
98 49 05 07 98 C9 83 C6 17 00 85 07 E9 CA 13 07
C0 02 63 8B E6 10 13 F7 F6 0D 13 06 50 04 63 1A
C7 08 D8 49 93 86 17 00 05 07 D8 C9 03 C7 17 00
63 06 07 10 13 06 C0 02 63 04 C7 10 D4 45 13 07
57 FD 13 77 D7 0F 85 06 D4 C5 25 E3 03 C7 27 00
93 86 27 00 75 C3 63 0D C7 0E 90 4D 13 07 07 FD
13 77 F7 0F 05 06 25 48 90 CD 63 78 E8 00 93 86
37 00 85 47 14 C1 3E 85 82 80 36 86 03 C7 16 00
85 06 93 08 C0 02 93 07 07 FD 93 F7 F7 0F 45 CF
63 0D 17 0B E3 73 F8 FE D8 41 85 47 93 06 26 00
3E 97 D8 C1 14 C1 3E 85 82 80 93 86 27 00 85 47
F5 B5 93 86 06 FD 93 F6 F6 0F 25 47 E3 75 D7 F4
D8 49 93 86 17 00 85 47 3E 97 D8 C9 C1 BD 90 41
93 87 16 00 05 06 90 C1 83 C6 16 00 9D FA BE 86
95 47 6D BD 81 47 85 06 55 BD 90 41 93 87 16 00
05 06 90 C1 03 C3 16 00 63 03 03 06 63 0D E3 04
90 45 13 07 03 FD 13 77 F7 0F A5 48 05 06 E3 F0
E8 EE 63 06 03 01 90 C5 89 06 85 47 41 B5 90 C5
DD B5 BE 86 91 47 9D BD BE 86 85 06 95 47 BD B5
BE 86 85 06 91 47 9D B5 99 47 8D B5 8D 47 B9 BD
8D 47 85 06 A1 BD 9D 47 91 BD 9D 47 85 06 B9 B5
99 47 85 06 A1 B5 BE 86 85 06 89 47 81 B5 BE 86
89 47 2D BD 19 71 CE D6 D2 D4 93 09 01 01 13 0A
01 03 A2 DC A6 DA CA D8 DA D0 DE CE E2 CC E6 CA
BE 84 3A 8B 86 DE D6 D2 2E 84 2E C6 AA 8C 32 8C
B6 8B D2 87 4E 89 4E 87 23 A0 07 00 23 20 07 00
91 07 94 08 11 07 E3 99 D7 FE 83 47 04 00 93 0A
C1 00 CD CF 0C 18 56 85 75 33 13 17 25 00 4E 97
B2 46 1C 43 83 C6 06 00 85 07 1C C3 E5 F6 22 C6
A2 9C 63 75 94 03 A2 87 13 06 C0 02 03 C7 07 00
B3 46 87 01 63 04 C7 00 23 80 D7 00 DA 97 E3 E7
97 FF 83 47 04 00 93 0A C1 00 91 CF 0C 18 56 85
95 33 13 17 25 00 4E 97 B2 46 1C 43 83 C6 06 00
85 07 1C C3 E5 F6 93 06 C0 02 63 7D 94 01 83 47
04 00 33 C7 77 01 63 84 D7 00 23 00 E4 00 5A 94
E3 67 94 FF 93 89 09 02 03 25 09 00 A6 85 11 09
01 26 AA 85 03 25 0A 00 11 0A DD 2C AA 84 E3 95
29 FF F6 50 66 54 D6 54 46 59 B6 59 26 5A 96 5A
06 5B F6 4B 66 4C D6 4C 09 61 82 80 A2 9C E3 64
94 F7 C9 B7 95 47 63 E4 A7 04 17 27 00 00 13 07
87 81 0A 05 3A 95 1C 41 BA 97 82 87 17 25 00 00
03 25 E5 C4 82 80 17 25 00 00 03 25 C5 C4 82 80
17 25 00 00 03 25 E5 C3 82 80 17 25 00 00 03 25
85 C1 82 80 17 25 00 00 03 25 A5 C0 82 80 01 45
82 80 13 F7 F5 0F 22 07 A1 81 85 67 7D 73 4D 8F
93 87 F7 F0 13 03 03 0F 33 76 F7 00 33 77 67 00
11 83 12 06 59 8E F5 78 0D 67 13 07 37 33 93 88
C8 CC 93 76 F5 00 B3 75 E6 00 11 81 33 76 16 01
92 06 C9 8E 09 82 8A 05 D1 8D 15 65 13 F6 36 03
6D 78 93 F6 C6 0C 13 08 A8 AA 13 DE 26 00 13 05
55 55 0A 06 B3 F6 A5 00 33 66 C6 01 B3 F5 05 01
85 81 86 06 93 7E 56 05 13 76 A6 0A 33 EE B6 00
86 0E 05 82 13 5E 8E 00 33 E6 CE 00 33 46 CE 00
06 06 17 1E 00 00 13 0E 8E 75 72 96 03 56 06 00
CD 8E A2 06 B1 8E 93 95 06 01 13 76 F6 0F 93 D6
85 01 22 06 55 8E B3 76 F6 00 33 76 66 00 11 82
92 06 D1 8E B3 F7 E6 00 B3 F6 16 01 89 82 8A 07
D5 8F 7D 8D B3 F7 07 01 85 83 06 05 5D 8D 82 80
93 F7 F5 0F A2 07 A1 81 05 67 7D 73 13 03 03 0F
13 07 F7 F0 CD 8F B3 F5 E7 00 B3 F7 67 00 91 83
92 05 DD 8D F5 78 8D 67 93 88 C8 CC 93 87 37 33
93 76 F5 00 13 78 05 0F 33 F6 F5 00 13 58 48 00
B3 F5 15 01 92 06 B3 E6 06 01 89 81 0A 06 4D 8E
13 FE 36 03 95 65 93 F6 C6 0C 6D 78 93 85 55 55
13 08 A8 AA 93 DE 26 00 0A 0E B3 76 B6 00 33 6E
DE 01 33 76 06 01 86 06 05 82 13 7F 5E 05 13 7E
AE 0A B3 EE C6 00 06 0F 13 5E 1E 00 93 DE 8E 00
33 6E CF 01 33 CE CE 01 55 8E 93 16 1E 00 17 1E
00 00 13 0E CE 66 F2 96 83 D6 06 00 22 06 21 81
35 8E 93 1E 06 01 93 F6 F6 0F 13 D6 8E 01 A2 06
D1 8E 33 F6 E6 00 B3 F6 66 00 91 82 12 06 55 8E
B3 76 F6 00 33 76 16 01 09 82 8A 06 D1 8E 33 F6
B6 00 B3 F6 06 01 06 06 85 82 D1 8E 13 F6 F6 0F
22 06 A1 82 55 8E B3 76 E6 00 B3 7E 66 00 93 DE
4E 00 13 76 F5 00 92 06 B3 E6 D6 01 11 81 12 06
49 8E B3 FE 16 01 33 F5 F6 00 93 DE 2E 00 93 76
36 03 0A 05 13 76 C6 0C 33 65 D5 01 09 82 8A 06
D1 8E 33 76 B5 00 33 75 05 01 13 FF 56 05 06 06
05 81 93 F6 A6 0A B3 6E A6 00 85 82 06 0F 33 6F
DF 00 93 D6 8E 00 B3 C6 E6 01 86 06 F2 96 83 D6
06 00 13 96 8E 00 35 8E 13 15 06 01 93 F6 F6 0F
13 56 85 01 A2 06 D1 8E 75 8F B3 F6 66 00 91 82
12 07 55 8F F9 8F 33 77 17 01 09 83 8A 07 D9 8F
33 F5 B7 00 B3 F7 07 01 85 83 06 05 5D 8D 82 80
93 F7 F5 0F A2 07 A1 81 05 67 FD 78 93 88 08 0F
13 07 F7 F0 CD 8F B3 F6 E7 00 B3 F7 17 01 91 83
92 06 DD 8E 75 78 8D 67 13 08 C8 CC 93 87 37 33
13 76 F5 00 93 75 05 0F 33 F3 F6 00 91 81 B3 F6
06 01 12 06 4D 8E 89 82 0A 03 33 63 D3 00 13 7E
36 03 95 66 13 76 C6 0C ED 75 93 86 56 55 93 85
A5 AA 93 5E 26 00 0A 0E 33 76 D3 00 33 6E DE 01
33 73 B3 00 06 06 13 53 13 00 13 7F 5E 05 13 7E
AE 0A B3 6E 66 00 06 0F 13 5E 1E 00 33 6E CF 01
93 DE 8E 00 B3 CE CE 01 33 6E 66 00 17 13 00 00
13 03 E3 4C 13 96 1E 00 1A 96 03 56 06 00 22 0E
13 5F 85 00 33 4E C6 01 93 1E 0E 01 13 76 F6 0F
13 DE 8E 01 22 06 33 66 C6 01 33 7E E6 00 33 76
16 01 11 82 12 0E 33 6E CE 00 33 76 FE 00 33 7E
0E 01 13 5E 2E 00 0A 06 33 66 C6 01 33 7E D6 00
6D 8E 05 82 06 0E 33 6E CE 00 13 76 FE 0F 22 06
13 5E 8E 00 33 66 C6 01 B3 7E E6 00 33 76 16 01
11 82 92 0E B3 EE CE 00 13 76 FF 00 13 7F 0F 0F
33 FE FE 00 13 5F 4F 00 B3 FE 0E 01 12 06 33 66
E6 01 93 DE 2E 00 0A 0E 33 6E DE 01 93 7E 36 03
13 76 C6 0C 13 5F 26 00 8A 0E 33 76 DE 00 B3 EE
EE 01 33 7E BE 00 06 06 13 5E 1E 00 93 FF 5E 05
93 FE AE 0A 33 6F C6 01 86 0F 93 DE 1E 00 13 5F
8F 00 B3 EE DF 01 B3 4E DF 01 33 6E C6 01 13 96
1E 00 1A 96 03 56 06 00 22 0E 93 5E 05 01 33 4E
C6 01 13 1F 0E 01 13 76 F6 0F 13 5E 8F 01 22 06
33 66 C6 01 33 7E E6 00 33 76 16 01 11 82 12 0E
33 6E CE 00 33 76 FE 00 33 7E 0E 01 13 5E 2E 00
0A 06 33 66 C6 01 33 7E D6 00 6D 8E 06 0E 05 82
33 66 CE 00 13 7E F6 0F 22 0E 21 82 33 6E CE 00
33 76 EE 00 33 7E 1E 01 13 5E 4E 00 12 06 33 66
C6 01 13 FE FE 00 93 FE 0E 0F 13 DF 4E 00 12 0E
B3 7E F6 00 33 76 06 01 33 6E EE 01 09 82 8A 0E
B3 EE CE 00 13 76 3E 03 13 7E CE 0C 13 5F 2E 00
0A 06 33 FE DE 00 33 66 E6 01 B3 FE BE 00 93 DE
1E 00 06 0E 93 7F 56 05 13 76 A6 0A 33 6F DE 01
86 0F 05 82 13 5F 8F 00 33 E6 CF 00 33 46 CF 00
06 06 1A 96 03 56 06 00 33 6E DE 01 22 0E 33 4E
C6 01 93 1E 0E 01 13 76 F6 0F 13 DE 8E 01 22 06
33 66 C6 01 33 7E E6 00 33 76 16 01 11 82 12 0E
33 6E CE 00 33 76 FE 00 33 7E 0E 01 13 5E 2E 00
0A 06 33 66 C6 01 33 7E D6 00 6D 8E 05 82 06 0E
33 6E CE 00 13 76 FE 0F 22 06 13 5E 8E 00 33 66
C6 01 B3 7E E6 00 33 7E 16 01 61 81 13 76 F5 00
13 5E 4E 00 92 0E 12 06 B3 EE CE 01 11 81 33 FE
FE 00 51 8D B3 FE 0E 01 13 76 35 03 93 DE 2E 00
13 75 C5 0C 0A 0E 33 6E DE 01 09 81 0A 06 49 8E
33 75 DE 00 33 7E BE 00 13 7F 56 05 06 05 13 5E
1E 00 13 76 A6 0A B3 6E C5 01 05 82 06 0F 33 6F
CF 00 13 D6 8E 00 33 46 E6 01 06 06 1A 96 03 56
06 00 13 95 8E 00 31 8D 13 13 05 01 13 76 F6 0F
13 55 83 01 22 06 49 8E 71 8F 33 76 16 01 11 82
12 07 51 8F F9 8F 33 77 07 01 09 83 8A 07 D9 8F
33 F5 D7 00 ED 8F 85 83 06 05 5D 8D 82 80 93 F7
F5 0F A2 07 A1 81 05 67 7D 73 13 03 03 0F 13 07
F7 F0 CD 8F B3 F5 E7 00 B3 F7 67 00 91 83 92 05
DD 8D F5 78 8D 67 93 88 C8 CC 93 87 37 33 93 76
F5 00 13 78 05 0F 33 F6 F5 00 13 58 48 00 B3 F5
15 01 92 06 B3 E6 06 01 89 81 0A 06 4D 8E 13 FE
36 03 95 65 93 F6 C6 0C 6D 78 93 85 55 55 13 08
A8 AA 93 DE 26 00 0A 0E B3 76 B6 00 33 6E DE 01
33 76 06 01 86 06 05 82 13 7F 5E 05 13 7E AE 0A
B3 EE C6 00 06 0F 13 5E 1E 00 93 DE 8E 00 33 6E
CF 01 33 CE CE 01 55 8E 93 16 1E 00 17 1E 00 00
13 0E EE 16 F2 96 83 D6 06 00 22 06 21 81 35 8E
93 1E 06 01 93 F6 F6 0F 13 D6 8E 01 A2 06 D1 8E
33 F6 E6 00 B3 F6 66 00 91 82 12 06 55 8E B3 76
F6 00 33 76 16 01 09 82 8A 06 D1 8E 33 F6 B6 00
B3 F6 06 01 06 06 85 82 D1 8E 13 F6 F6 0F 22 06
A1 82 55 8E B3 76 E6 00 B3 7E 66 00 93 DE 4E 00
13 76 F5 00 92 06 13 75 05 0F B3 E6 D6 01 11 81
12 06 49 8E B3 FE 16 01 33 F5 F6 00 93 DE 2E 00
93 76 36 03 0A 05 13 76 C6 0C 33 65 D5 01 09 82
8A 06 D1 8E 33 76 B5 00 33 75 05 01 13 FF 56 05
06 06 05 81 93 F6 A6 0A B3 6E A6 00 85 82 06 0F
33 6F DF 00 93 D6 8E 00 B3 C6 E6 01 86 06 F2 96
83 D6 06 00 13 96 8E 00 35 8E 13 15 06 01 93 F6
F6 0F 13 56 85 01 A2 06 D1 8E 75 8F B3 F6 66 00
91 82 12 07 55 8F F9 8F 33 77 17 01 09 83 8A 07
D9 8F 33 F5 B7 00 B3 F7 07 01 85 83 06 05 5D 8D
82 80 01 45 82 80 B7 07 D9 00 8D 07 37 07 00 20
1C C3 82 80 B7 02 00 30 83 A5 42 00 03 A5 02 00
03 A3 42 00 E3 98 65 FE 82 80 B7 02 00 30 83 A7
42 00 03 A7 02 00 03 A3 42 00 E3 98 67 FE 97 16
00 00 23 AA E6 44 17 17 00 00 23 28 F7 44 82 80
B7 02 00 30 83 A7 42 00 03 A7 02 00 03 A3 42 00
E3 98 67 FE 97 16 00 00 23 A3 E6 42 17 17 00 00
23 21 F7 42 82 80 97 16 00 00 93 86 46 41 17 17
00 00 13 07 47 41 9C 42 08 43 CC 42 58 43 33 85
A7 40 B3 B7 A7 00 99 8D 9D 8D 82 80 B7 47 E6 55
93 87 97 B8 33 35 F5 02 5D 81 82 80 B7 07 D9 00
8D 07 37 07 00 20 1C C3 85 47 23 00 F5 00 82 80
23 00 05 00 82 80 1D 71 A2 CE A6 CC 13 F8 07 04
97 1F 00 00 93 8F 6F EC 63 06 08 00 97 1F 00 00
93 8F 2F EE 93 F3 07 01 63 96 03 0A 13 F4 17 00
93 0E F4 FF 93 FE 0E FF 93 8E 0E 03 13 F8 27 00
93 F2 07 02 63 06 08 08 63 C1 05 1A 13 F8 47 00
63 1E 08 16 A1 8B 81 44 81 C7 FD 16 93 04 00 02
63 8C 02 00 C1 47 63 02 F6 1A 93 07 86 FF 93 B7
17 00 9D 8E 93 02 00 02 63 9B 05 10 93 07 00 03
23 06 F1 00 01 4F 05 48 93 08 C1 00 42 8E 63 53
E8 00 3A 8E B3 86 C6 41 21 E4 33 03 D5 00 AA 87
93 05 00 02 63 5D D0 02 85 07 A3 8F B7 FE E3 9D
67 FE 3E 85 63 91 04 10 63 88 02 00 A1 46 63 08
D6 16 C1 46 63 08 D6 10 B3 36 70 00 F9 16 99 A0
81 44 79 B7 F9 9B 41 44 93 0E 00 02 85 B7 FD 16
81 C4 23 00 95 00 05 05 63 88 02 00 A1 47 63 02
F6 12 C1 47 63 01 F6 0E 63 9E 03 00 33 06 D5 00
AA 87 63 52 D0 14 85 07 A3 8F D7 FF E3 9D C7 FE
3E 85 FD 56 AA 87 33 03 C5 01 93 05 00 03 63 51
E8 02 85 07 33 06 F3 40 A3 8F B7 FE E3 4B C8 FE
81 47 63 55 E8 00 B3 07 0E 41 FD 17 85 07 3E 95
B3 87 E8 01 93 85 F8 FF 2A 87 03 C6 07 00 FD 17
05 07 A3 0F C7 FE E3 9A F5 FE B3 07 E5 01 93 85
17 00 2E 85 63 5E D0 00 13 87 16 00 3E 97 13 06
00 02 23 00 C5 00 05 05 E3 1D A7 FE 33 85 B6 00
76 44 E6 44 25 61 82 80 FD 16 93 04 D0 02 01 48
93 08 C1 00 B3 F7 C5 02 42 8F 05 08 33 8E 08 01
2E 83 FE 97 83 C7 07 00 B3 D5 C5 02 A3 0F FE FE
E3 72 C3 FE E1 BD 23 80 97 00 13 85 17 00 63 90
02 06 F9 56 E3 88 03 F4 FD 56 A9 B7 FD 16 93 04
B0 02 79 B5 FD 56 13 06 00 03 93 07 80 07 23 00
C5 00 A3 00 F5 00 09 05 01 BF B3 05 B0 40 E3 8D
02 F8 C1 47 63 03 F6 04 A1 47 63 04 F6 02 FD 16
93 04 D0 02 93 02 00 02 59 B7 F9 16 93 02 00 02
A5 B5 93 07 00 03 23 00 F5 00 05 05 F1 BD FD 56
F1 B5 F9 16 93 04 D0 02 93 02 00 02 8D B7 93 07
00 03 23 00 F5 00 05 05 69 B7 F5 16 93 04 D0 02
93 02 00 02 A9 B7 FD 16 F1 B5 B7 07 00 20 C8 43
05 89 82 80 37 07 00 20 11 07 1C 43 85 8B F5 FF
B7 07 00 20 C8 C7 82 80 83 46 05 00 99 CE 37 07
00 20 37 06 00 20 11 07 31 06 05 05 1C 43 85 8B
F5 FF 14 C2 83 46 05 00 ED FA 82 80 37 07 00 20
11 07 1C 43 85 8B F5 FF B7 07 00 20 C8 C7 82 80
13 01 01 B8 23 28 21 45 23 2E 11 44 23 26 31 45
23 22 B1 46 23 24 C1 46 23 26 D1 46 23 28 E1 46
23 2A F1 46 23 2C 01 47 23 2E 11 47 83 47 05 00
13 09 41 46 4A CA 63 8C 07 60 93 09 01 03 23 2C
81 44 23 2A 91 44 23 24 41 45 23 22 51 45 23 20
61 45 23 2E 71 43 2A 83 23 2C 81 43 4E 85 13 0A
50 02 C1 44 17 14 00 00 13 04 64 EA A5 4B 13 0B
E0 02 93 0A C0 04 63 8D 47 05 23 00 F5 00 83 47
13 00 05 05 05 03 E5 FB 03 24 81 45 83 24 41 45
03 2A 81 44 83 2A 41 44 03 2B 01 44 83 2B C1 43
03 2C 81 43 23 00 05 00 03 46 01 03 63 0A 06 5A
37 07 00 20 B7 05 00 20 11 07 B1 05 CE 86 1C 43
85 8B F5 FF 90 C1 03 C6 16 00 61 CE 85 06 C5 BF
81 47 03 46 13 00 13 08 13 00 13 07 06 FE 13 77
F7 0F 63 E7 E4 00 0A 07 22 97 18 43 22 97 02 87
13 07 06 FD 13 77 F7 0F 63 F4 EB 0E 13 07 A0 02
FD 56 63 02 E6 10 7D 57 63 0A 66 0B 93 75 F6 0D
63 98 55 07 32 83 03 46 18 00 93 08 70 03 13 0C
18 00 93 05 F6 FB 93 F5 F5 0F 63 EF B8 02 97 18
00 00 93 88 08 E2 8A 05 C6 95 8C 41 C6 95 82 85
93 E7 17 00 42 83 71 B7 93 E7 07 01 42 83 51 B7
93 E7 47 00 42 83 B5 BF 93 E7 07 02 42 83 95 BF
93 E7 87 00 42 83 B5 B7 62 88 93 07 50 02 63 03
F6 20 23 00 F5 00 83 47 08 00 05 05 91 D7 ED AA
93 05 F6 FB 93 F5 F5 0F 93 08 70 03 E3 EF B8 FC
97 18 00 00 93 88 E8 E9 8A 05 C6 95 8C 41 C6 95
82 85 83 20 C1 45 B3 86 36 41 03 29 01 45 83 29
C1 44 13 85 16 00 13 01 01 48 82 80 03 46 18 00
25 43 93 05 18 00 13 07 06 FD 13 77 F7 0F 63 70
E3 16 13 07 A0 02 63 04 E6 18 2E 88 01 47 3D B7
81 46 A5 45 13 97 26 00 36 97 05 08 06 07 32 97
03 46 08 00 93 06 07 FD 13 07 06 FD 13 77 F7 0F
E3 F2 E5 FE 09 B7 83 26 09 00 03 46 23 00 13 08
23 00 63 C4 06 00 11 09 FD B5 B3 06 D0 40 93 E7
07 01 11 09 CD B5 93 E7 07 04 41 46 83 25 09 00
11 09 15 3E 83 47 1C 00 13 03 1C 00 E3 9D 07 E2
A1 B5 42 8C 29 46 DD B7 62 88 C1 8B 93 05 49 00
13 03 18 00 63 86 07 14 83 27 09 00 13 06 15 00
85 48 23 00 F5 00 13 07 00 02 36 95 B2 87 63 D7
D8 46 85 07 A3 8F E7 FE E3 9D A7 FE FD 16 33 05
D6 00 83 47 18 00 2E 89 E3 97 07 DE F5 BB 62 88
03 26 09 00 11 09 63 0F 06 0E 83 45 06 00 C1 8B
63 80 05 42 B3 08 E6 00 32 87 63 07 17 01 83 45
17 00 05 07 FD F9 BA 88 B3 88 C8 40 63 88 07 10
63 5E 10 01 B3 05 16 01 AA 87 03 47 06 00 05 06
85 07 A3 8F E7 FE E3 1A B6 FE 46 95 33 87 16 41
2A 97 13 03 18 00 AA 87 13 06 00 02 63 DA D8 00
85 07 A3 8F C7 FE E3 9D E7 FE AA 96 33 85 16 41
83 47 18 00 E3 99 07 D6 41 B3 62 88 7D 56 63 8F
C6 06 83 25 09 00 41 46 42 C6 B1 34 32 48 11 09
83 47 18 00 13 03 18 00 E3 97 07 D4 B1 BB 81 48
13 97 28 00 46 97 85 05 06 07 32 97 03 C6 05 00
93 08 07 FD 13 07 06 FD 13 77 F7 0F E3 72 E3 FE
13 C7 F8 FF 7D 87 2E 88 33 F7 E8 00 45 BB 03 27
09 00 03 46 28 00 11 09 93 45 F7 FF FD 85 6D 8F
09 08 69 BB 83 47 08 00 23 00 F5 00 83 47 18 00
05 05 13 03 18 00 E3 98 07 CE FD B9 93 E7 17 00
A1 46 41 B7 C1 8B 17 16 00 00 13 06 06 8F 19 B7
85 47 63 D4 D7 30 13 87 F6 FF 2A 97 AA 87 13 06
00 02 85 07 A3 8F C7 FE E3 1D F7 FE 83 27 09 00
7D 15 36 95 23 00 F5 00 05 05 65 BD 63 DD D8 2C
33 87 16 41 2A 97 AA 87 93 05 00 02 85 07 A3 8F
B7 FE E3 9D E7 FE AA 96 33 85 16 41 93 86 F8 FF
C1 BD 13 06 C0 06 93 E7 27 00 E3 05 C3 E4 83 25
09 00 29 46 11 09 35 B5 13 07 C0 06 63 04 E3 26
03 2E 09 00 11 09 03 46 0E 00 63 03 06 22 01 48
81 48 05 47 93 05 30 06 63 DE C5 1C B7 85 EB 51
93 85 F5 51 B3 35 B6 02 13 0F 40 06 17 03 00 00
13 03 A3 7F B7 DE CC CC 93 8E DE CC 0A 97 95 81
33 8F E5 03 9A 95 83 CF 05 00 B3 85 28 00 89 08
23 8C F5 01 B3 05 E6 41 33 B6 D5 03 0D 82 B3 0E
C3 00 03 CF 0E 00 93 1E 26 00 76 96 06 06 23 0C
E7 01 33 86 C5 40 33 07 C3 00 83 45 07 00 33 86
28 00 05 08 23 0C B6 00 11 46 13 87 18 00 63 09
C8 02 33 06 0E 01 03 46 06 00 B3 05 27 00 93 08
E0 02 23 8C 15 01 93 08 17 00 09 07 25 F6 13 06
00 03 8A 98 23 8C C8 00 05 08 11 46 E3 1B C8 FC
C1 8B 9D E3 63 50 D7 20 33 86 E6 40 2A 96 AA 87
93 05 00 02 85 07 A3 8F B7 FE E3 9D C7 FE AA 96
33 85 E6 40 93 06 F7 FF 63 5D E0 00 3C 08 B3 05
E5 00 03 C6 07 00 05 05 85 07 A3 0F C5 FE E3 1A
B5 FE E3 51 D7 D2 B3 87 E6 40 AA 97 13 07 00 02
05 05 A3 0F E5 FE E3 1D F5 FE 29 B3 13 07 C0 06
93 E7 07 04 E3 1E E3 EC 83 2E 09 00 17 03 00 00
13 03 23 72 11 09 81 48 01 46 19 4F 93 0F A0 03
29 A0 96 95 23 84 F5 01 0D 06 33 87 1E 01 03 47
07 00 93 02 01 01 85 08 93 55 47 00 9A 95 03 CE
05 00 3D 8B 1A 97 83 45 07 00 33 07 56 00 23 04
C7 01 13 0E 16 00 33 07 5E 00 23 04 B7 00 93 05
26 00 E3 90 E8 FD C1 8B 95 E3 B3 87 B6 40 AA 97
2A 87 13 06 00 02 63 D9 D5 12 05 07 A3 0F C7 FE
E3 1D F7 FE AA 96 33 85 B6 40 F2 86 3C 08 33 06
B5 00 03 C7 07 00 05 05 85 07 A3 0F E5 FE E3 1A
C5 FE 63 DF D5 00 B3 87 B6 40 B3 06 F6 00 13 07
00 02 05 05 A3 0F E5 FE E3 9D A6 FE 33 05 F6 00
83 47 28 00 13 03 28 00 E3 9F 07 A6 71 B4 42 8C
21 46 2D B1 A5 45 17 03 00 00 13 03 03 63 E3 DC
C5 E6 B7 D5 CC CC 93 85 D5 CC B3 35 B6 02 B3 8E
28 00 BA 88 13 D7 35 00 B3 05 E3 00 03 CF 05 00
93 15 27 00 2E 97 06 07 23 8C EE 01 19 8E A1 B5
13 07 00 03 23 0C E1 00 05 47 3A 88 99 BD 93 09
01 03 4E 85 23 00 05 00 03 46 01 03 E3 1A 06 A4
83 20 C1 45 03 29 01 45 83 29 C1 44 01 45 13 01
01 48 82 80 83 2E 09 00 17 03 00 00 13 03 E3 5B
11 09 D1 B5 93 E7 27 00 42 8C 95 BB 42 8C 49 B3
42 8C 61 BE 93 E7 07 04 42 8C 9D BB 93 E7 07 04
42 8C 41 46 61 B6 FD 16 21 B9 83 27 09 00 05 05
2E 89 A3 0F F5 FE 83 47 18 00 E3 9E 07 9A E9 B2
81 48 E3 9D 07 C0 13 03 18 00 E3 43 D0 D0 83 47
18 00 0D B9 FD 16 0D B5 FD 16 CD B5 32 85 55 B6
@800027B8
36 6B 20 70 65 72 66 6F 72 6D 61 6E 63 65 20 72
75 6E 20 70 61 72 61 6D 65 74 65 72 73 20 66 6F
72 20 63 6F 72 65 6D 61 72 6B 2E 0A 00 00 00 00
36 6B 20 76 61 6C 69 64 61 74 69 6F 6E 20 72 75
6E 20 70 61 72 61 6D 65 74 65 72 73 20 66 6F 72
20 63 6F 72 65 6D 61 72 6B 2E 0A 00 50 72 6F 66
69 6C 65 20 67 65 6E 65 72 61 74 69 6F 6E 20 72
75 6E 20 70 61 72 61 6D 65 74 65 72 73 20 66 6F
72 20 63 6F 72 65 6D 61 72 6B 2E 0A 00 00 00 00
32 4B 20 70 65 72 66 6F 72 6D 61 6E 63 65 20 72
75 6E 20 70 61 72 61 6D 65 74 65 72 73 20 66 6F
72 20 63 6F 72 65 6D 61 72 6B 2E 0A 00 00 00 00
32 4B 20 76 61 6C 69 64 61 74 69 6F 6E 20 72 75
6E 20 70 61 72 61 6D 65 74 65 72 73 20 66 6F 72
20 63 6F 72 65 6D 61 72 6B 2E 0A 00 5B 25 75 5D
45 52 52 4F 52 21 20 6C 69 73 74 20 63 72 63 20
30 78 25 30 34 78 20 2D 20 73 68 6F 75 6C 64 20
62 65 20 30 78 25 30 34 78 0A 00 00 5B 25 75 5D
45 52 52 4F 52 21 20 6D 61 74 72 69 78 20 63 72
63 20 30 78 25 30 34 78 20 2D 20 73 68 6F 75 6C
64 20 62 65 20 30 78 25 30 34 78 0A 00 00 00 00
5B 25 75 5D 45 52 52 4F 52 21 20 73 74 61 74 65
20 63 72 63 20 30 78 25 30 34 78 20 2D 20 73 68
6F 75 6C 64 20 62 65 20 30 78 25 30 34 78 0A 00
43 6F 72 65 4D 61 72 6B 20 53 69 7A 65 20 20 20
20 3A 20 25 6C 75 0A 00 54 6F 74 61 6C 20 74 69
63 6B 73 20 20 20 20 20 20 3A 20 25 6C 75 0A 00
54 6F 74 61 6C 20 74 69 6D 65 20 28 73 65 63 73
29 3A 20 25 64 0A 00 00 49 74 65 72 61 74 69 6F
6E 73 2F 53 65 63 20 20 20 3A 20 25 64 0A 00 00
45 52 52 4F 52 21 20 4D 75 73 74 20 65 78 65 63
75 74 65 20 66 6F 72 20 61 74 20 6C 65 61 73 74
20 31 30 20 73 65 63 73 20 66 6F 72 20 61 20 76
61 6C 69 64 20 72 65 73 75 6C 74 21 0A 00 00 00
49 74 65 72 61 74 69 6F 6E 73 20 20 20 20 20 20
20 3A 20 25 6C 75 0A 00 47 43 43 31 35 2E 31 2E
30 00 00 00 43 6F 6D 70 69 6C 65 72 20 76 65 72
73 69 6F 6E 20 3A 20 25 73 0A 00 00 2D 4F 32 20
2D 6D 63 6D 6F 64 65 6C 3D 6D 65 64 61 6E 79 20
2D 73 74 64 3D 67 6E 75 39 39 20 2D 66 6E 6F 2D
63 6F 6D 6D 6F 6E 20 2D 66 6E 6F 2D 62 75 69 6C
74 69 6E 20 2D 66 66 75 6E 63 74 69 6F 6E 2D 73
65 63 74 69 6F 6E 73 20 2D 44 50 45 52 46 4F 52
4D 41 4E 43 45 5F 52 55 4E 3D 31 20 20 2D 6E 6F
73 74 64 6C 69 62 20 2D 6E 6F 73 74 61 72 74 66
69 6C 65 73 20 2D 73 74 61 74 69 63 20 2D 54 20
72 76 33 32 69 6D 63 2D 62 61 72 65 6D 65 74 61
6C 2F 6C 69 6E 6B 2E 6C 64 20 2D 6C 6D 20 2D 6C
67 63 63 00 43 6F 6D 70 69 6C 65 72 20 66 6C 61
67 73 20 20 20 3A 20 25 73 0A 00 00 53 54 41 43
4B 00 00 00 4D 65 6D 6F 72 79 20 6C 6F 63 61 74
69 6F 6E 20 20 3A 20 25 73 0A 00 00 73 65 65 64
63 72 63 20 20 20 20 20 20 20 20 20 20 3A 20 30
78 25 30 34 78 0A 00 00 5B 25 64 5D 63 72 63 6C
69 73 74 20 20 20 20 20 20 20 3A 20 30 78 25 30
34 78 0A 00 5B 25 64 5D 63 72 63 6D 61 74 72 69
78 20 20 20 20 20 3A 20 30 78 25 30 34 78 0A 00
5B 25 64 5D 63 72 63 73 74 61 74 65 20 20 20 20
20 20 3A 20 30 78 25 30 34 78 0A 00 5B 25 64 5D
63 72 63 66 69 6E 61 6C 20 20 20 20 20 20 3A 20
30 78 25 30 34 78 0A 00 43 6F 72 72 65 63 74 20
6F 70 65 72 61 74 69 6F 6E 20 76 61 6C 69 64 61
74 65 64 2E 20 53 65 65 20 52 45 41 44 4D 45 2E
6D 64 20 66 6F 72 20 72 75 6E 20 61 6E 64 20 72
65 70 6F 72 74 69 6E 67 20 72 75 6C 65 73 2E 0A
00 00 00 00 43 61 6E 6E 6F 74 20 76 61 6C 69 64
61 74 65 20 6F 70 65 72 61 74 69 6F 6E 20 66 6F
72 20 74 68 65 73 65 20 73 65 65 64 20 76 61 6C
75 65 73 2C 20 70 6C 65 61 73 65 20 63 6F 6D 70
61 72 65 20 77 69 74 68 20 72 65 73 75 6C 74 73
20 6F 6E 20 61 20 6B 6E 6F 77 6E 20 70 6C 61 74
66 6F 72 6D 2E 0A 00 00 45 72 72 6F 72 73 20 64
65 74 65 63 74 65 64 0A 00 00 00 00 53 74 61 74
69 63 00 00 48 65 61 70 00 00 00 00 53 74 61 63
6B 00 00 00 54 30 2E 33 65 2D 31 46 00 00 00 00
2D 54 2E 54 2B 2B 54 71 00 00 00 00 31 54 33 2E
34 65 34 7A 00 00 00 00 33 34 2E 30 65 2D 54 5E
00 00 00 00 35 2E 35 30 30 65 2B 33 00 00 00 00
2D 2E 31 32 33 65 2D 32 00 00 00 00 2D 38 37 65
2B 38 33 32 00 00 00 00 2B 30 2E 36 65 2D 31 32
00 00 00 00 33 35 2E 35 34 34 30 30 00 00 00 00
2E 31 32 33 34 35 30 30 00 00 00 00 2D 31 31 30
2E 37 30 30 00 00 00 00 2B 30 2E 36 34 34 30 30
00 00 00 00 35 30 31 32 00 00 00 00 31 32 33 34
00 00 00 00 2D 38 37 34 00 00 00 00 2B 31 32 32
00 00 00 00 30 31 32 33 34 35 36 37 38 39 61 62
63 64 65 66 67 68 69 6A 6B 6C 6D 6E 6F 70 71 72
73 74 75 76 77 78 79 7A 00 00 00 00 30 31 32 33
34 35 36 37 38 39 41 42 43 44 45 46 47 48 49 4A
4B 4C 4D 4E 4F 50 51 52 53 54 55 56 57 58 59 5A
00 00 00 00 3C 4E 55 4C 4C 3E 00 00 B0 D4 40 33
79 6A 14 E7 C1 E3 00 00 52 BE 99 11 08 56 D7 1F
47 07 00 00 47 5E BF 39 A4 E5 3A 8E 84 8D 00 00
EC 2C 00 80 F4 2C 00 80 FC 2C 00 80 04 2D 00 80
BC 2C 00 80 C8 2C 00 80 D4 2C 00 80 E0 2C 00 80
8C 2C 00 80 98 2C 00 80 A4 2C 00 80 B0 2C 00 80
5C 2C 00 80 68 2C 00 80 74 2C 00 80 80 2C 00 80
2C E8 FF FF 04 E8 FF FF 0E E8 FF FF 18 E8 FF FF
22 E8 FF FF FA E7 FF FF 00 00 05 80 0F 80 0A 00
1B 80 1E 00 14 00 11 80 33 80 36 00 3C 00 39 80
28 00 2D 80 27 80 22 00 63 80 66 00 6C 00 69 80
78 00 7D 80 77 80 72 00 50 00 55 80 5F 80 5A 00
4B 80 4E 00 44 00 41 80 C3 80 C6 00 CC 00 C9 80
D8 00 DD 80 D7 80 D2 00 F0 00 F5 80 FF 80 FA 00
EB 80 EE 00 E4 00 E1 80 A0 00 A5 80 AF 80 AA 00
BB 80 BE 00 B4 00 B1 80 93 80 96 00 9C 00 99 80
88 00 8D 80 87 80 82 00 83 81 86 01 8C 01 89 81
98 01 9D 81 97 81 92 01 B0 01 B5 81 BF 81 BA 01
AB 81 AE 01 A4 01 A1 81 E0 01 E5 81 EF 81 EA 01
FB 81 FE 01 F4 01 F1 81 D3 81 D6 01 DC 01 D9 81
C8 01 CD 81 C7 81 C2 01 40 01 45 81 4F 81 4A 01
5B 81 5E 01 54 01 51 81 73 81 76 01 7C 01 79 81
68 01 6D 81 67 81 62 01 23 81 26 01 2C 01 29 81
38 01 3D 81 37 81 32 01 10 01 15 81 1F 81 1A 01
0B 81 0E 01 04 01 01 81 03 83 06 03 0C 03 09 83
18 03 1D 83 17 83 12 03 30 03 35 83 3F 83 3A 03
2B 83 2E 03 24 03 21 83 60 03 65 83 6F 83 6A 03
7B 83 7E 03 74 03 71 83 53 83 56 03 5C 03 59 83
48 03 4D 83 47 83 42 03 C0 03 C5 83 CF 83 CA 03
DB 83 DE 03 D4 03 D1 83 F3 83 F6 03 FC 03 F9 83
E8 03 ED 83 E7 83 E2 03 A3 83 A6 03 AC 03 A9 83
B8 03 BD 83 B7 83 B2 03 90 03 95 83 9F 83 9A 03
8B 83 8E 03 84 03 81 83 80 02 85 82 8F 82 8A 02
9B 82 9E 02 94 02 91 82 B3 82 B6 02 BC 02 B9 82
A8 02 AD 82 A7 82 A2 02 E3 82 E6 02 EC 02 E9 82
F8 02 FD 82 F7 82 F2 02 D0 02 D5 82 DF 82 DA 02
CB 82 CE 02 C4 02 C1 82 43 82 46 02 4C 02 49 82
58 02 5D 82 57 82 52 02 70 02 75 82 7F 82 7A 02
6B 82 6E 02 64 02 61 82 20 02 25 82 2F 82 2A 02
3B 82 3E 02 34 02 31 82 13 82 16 02 1C 02 19 82
08 02 0D 82 07 82 02 02 56 F2 FF FF E6 F1 FF FF
E6 F1 FF FF 4E F2 FF FF E6 F1 FF FF E6 F1 FF FF
E6 F1 FF FF E6 F1 FF FF E6 F1 FF FF E6 F1 FF FF
E6 F1 FF FF 46 F2 FF FF E6 F1 FF FF 3E F2 FF FF
E6 F1 FF FF E6 F1 FF FF 36 F2 FF FF DE F5 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF D8 F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF BA F4 FF FF
1A F2 FF FF FA F2 FF FF A4 F4 FF FF 1A F2 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF A4 F4 FF FF
1A F2 FF FF 1A F2 FF FF 1A F2 FF FF 1A F2 FF FF
1A F2 FF FF B2 F6 FF FF BC F3 FF FF 1A F2 FF FF
1A F2 FF FF 40 F3 FF FF 1A F2 FF FF F6 F2 FF FF
1A F2 FF FF 1A F2 FF FF DC F2 FF FF 66 F6 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 6E F6 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 5E F6 FF FF
3C F1 FF FF 1C F2 FF FF 56 F6 FF FF 3C F1 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 56 F6 FF FF
3C F1 FF FF 3C F1 FF FF 3C F1 FF FF 3C F1 FF FF
3C F1 FF FF D0 F5 FF FF DE F2 FF FF 3C F1 FF FF
3C F1 FF FF 62 F2 FF FF 3C F1 FF FF 14 F2 FF FF
3C F1 FF FF 3C F1 FF FF 62 F6 FF FF
@800031E4
44 2C 00 80 4C 2C 00 80 54 2C 00 80 01 00 00 00
D0 07 00 00 66 00 00 00
