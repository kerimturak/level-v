/*
Copyright (c) 2025 Kerim TURAK

Permission is granted to use, copy, modify, and distribute this software for any purpose,
with or without fee, provided that the above notice appears in all copies.

THE SOFTWARE IS PROVIDED "AS IS" WITHOUT ANY WARRANTY OF ANY KIND.

Description:
  Word-based (32-bit) RAM with cache line burst support.
  
  Features:
    - 32-bit word organization (standard .mem file compatible)
    - Cache line width read/write (128-bit default)
    - UART programming interface via separate module
    - Configurable depth and timing
  
  Memory Organization:
    - Words are 32-bit aligned
    - Cache lines span WORDS_PER_LINE consecutive words
    - Byte strobes enable fine-grained writes
*/
`timescale 1ns / 1ps

module wrapper_ram
  import ceres_param::*;
#(
    // Memory Configuration
    parameter int unsigned WORD_WIDTH       = 32,
    parameter int unsigned RAM_DEPTH        = 32768,
    parameter int unsigned CACHE_LINE_WIDTH = BLK_SIZE,

    // Programming Configuration  
    parameter int unsigned                              CPU_CLK          = ceres_param::CPU_CLK,
    parameter int unsigned                              PROG_BAUD_RATE   = ceres_param::PROG_BAUD_RATE,
    parameter logic        [8*PROGRAM_SEQUENCE_LEN-1:0] PROGRAM_SEQUENCE = ceres_param::PROGRAM_SEQUENCE
) (
    input logic clk_i,
    input logic rst_ni,

    // Memory Interface (cache line width)
    input  logic [ $clog2(RAM_DEPTH)-1:0] addr_i,
    input  logic [  CACHE_LINE_WIDTH-1:0] wdata_i,
    input  logic [CACHE_LINE_WIDTH/8-1:0] wstrb_i,
    output logic [  CACHE_LINE_WIDTH-1:0] rdata_o,
    input  logic                          rd_en_i,

    // Programming Interface
    input  logic ram_prog_rx_i,
    output logic system_reset_o,
    output logic prog_mode_led_o
);

  // ==========================================================================
  // Derived Parameters
  // ==========================================================================
  localparam int WORDS_PER_LINE = CACHE_LINE_WIDTH / WORD_WIDTH;
  localparam int BYTES_PER_WORD = WORD_WIDTH / 8;
  localparam int LINE_ADDR_BITS = $clog2(WORDS_PER_LINE);

  // ==========================================================================
  // Memory Array - Separate BRAMs for each word position
  // ==========================================================================
  // Split into individual BRAMs for proper inference
  (* ram_style = "block" *)logic [                      WORD_WIDTH-1:0] ram0         [RAM_DEPTH/WORDS_PER_LINE-1:0];
  (* ram_style = "block" *)logic [                      WORD_WIDTH-1:0] ram1         [RAM_DEPTH/WORDS_PER_LINE-1:0];
  (* ram_style = "block" *)logic [                      WORD_WIDTH-1:0] ram2         [RAM_DEPTH/WORDS_PER_LINE-1:0];
  (* ram_style = "block" *)logic [                      WORD_WIDTH-1:0] ram3         [RAM_DEPTH/WORDS_PER_LINE-1:0];

  // ==========================================================================
  // Internal Signals
  // ==========================================================================

  // Address calculation
  logic [$clog2(RAM_DEPTH/WORDS_PER_LINE)-1:0] word_addr;

  // Read data registers - separate for each BRAM to enable proper output register inference
  logic [                      WORD_WIDTH-1:0] rdata_q0;
  logic [                      WORD_WIDTH-1:0] rdata_q1;
  logic [                      WORD_WIDTH-1:0] rdata_q2;
  logic [                      WORD_WIDTH-1:0] rdata_q3;

  // Programming interface
  logic [                                31:0] prog_addr;
  logic [                                31:0] prog_data;
  logic                                        prog_valid;
  logic                                        prog_mode;
  logic                                        prog_sys_rst;

  // ==========================================================================
  // Memory Initialization
  // ==========================================================================
  localparam int INIT_FILE_LEN = 256;
  reg     [8*INIT_FILE_LEN-1:0] init_file = {INIT_FILE_LEN{8'h00}};
  integer                       fd = 0;
  logic   [     WORD_WIDTH-1:0] temp_ram                           [0:RAM_DEPTH-1];

  initial begin
`ifndef SYNTHESIS
    if ($value$plusargs("INIT_FILE=%s", init_file)) begin
      fd = $fopen(init_file, "r");
      if (fd == 0) begin
        $display("[ERROR] Cannot open memory file: %s", init_file);
        $finish;
      end
      $fclose(fd);
      $readmemh(init_file, temp_ram, 0, RAM_DEPTH - 1);
      // Distribute to separate BRAMs
      for (int i = 0; i < RAM_DEPTH; i += 4) begin
        ram0[i/4] = temp_ram[i];
        ram1[i/4] = temp_ram[i+1];
        ram2[i/4] = temp_ram[i+2];
        ram3[i/4] = temp_ram[i+3];
      end
`ifdef LOG_RAM
      $display("[INFO] Memory loaded successfully.");
`endif
    end else begin
`ifdef LOG_RAM
      $display("[INFO] No INIT_FILE -> RAM initialized to zero");
`endif
    end
`else
    // During synthesis, initialize to zero (BRAM will be initialized via .coe or programming interface)
    for (int i = 0; i < RAM_DEPTH / WORDS_PER_LINE; i++) begin
      ram0[i] = '0;
      ram1[i] = '0;
      ram2[i] = '0;
      ram3[i] = '0;
    end
`endif
  end

  // ==========================================================================
  // Address Calculation
  // ==========================================================================
  assign word_addr = addr_i[$clog2(RAM_DEPTH)-1:LINE_ADDR_BITS];

  // ==========================================================================
  // Read/Write Logic - BRAM-Friendly Template (UG901 Style)
  // ==========================================================================
  // Simplified to match Vivado BRAM inference patterns:
  // - Separate write enable and read enable
  // - No complex conditional logic in clocked block
  // - Write-first behavior through explicit output assignment

  // Write enable signals for each bank
  logic we0, we1, we2, we3;
  logic [$clog2(RAM_DEPTH/WORDS_PER_LINE)-1:0] wr_addr;
  logic [WORD_WIDTH-1:0] wr_data0, wr_data1, wr_data2, wr_data3;

  // Write enable and data muxing
  always_comb begin
    if (prog_mode && prog_valid) begin
      // Programming mode: write to specific bank based on address[1:0]
      wr_addr = prog_addr[$clog2(RAM_DEPTH)-1:LINE_ADDR_BITS];
      we0 = (prog_addr[LINE_ADDR_BITS-1:0] == 2'd0);
      we1 = (prog_addr[LINE_ADDR_BITS-1:0] == 2'd1);
      we2 = (prog_addr[LINE_ADDR_BITS-1:0] == 2'd2);
      we3 = (prog_addr[LINE_ADDR_BITS-1:0] == 2'd3);
      wr_data0 = prog_data;
      wr_data1 = prog_data;
      wr_data2 = prog_data;
      wr_data3 = prog_data;
    end else begin
      // Normal mode: write based on byte strobes
      wr_addr = word_addr;
      we0 = |wstrb_i[0*BYTES_PER_WORD+:BYTES_PER_WORD];
      we1 = |wstrb_i[1*BYTES_PER_WORD+:BYTES_PER_WORD];
      we2 = |wstrb_i[2*BYTES_PER_WORD+:BYTES_PER_WORD];
      we3 = |wstrb_i[3*BYTES_PER_WORD+:BYTES_PER_WORD];
      wr_data0 = wdata_i[0*WORD_WIDTH+:WORD_WIDTH];
      wr_data1 = wdata_i[1*WORD_WIDTH+:WORD_WIDTH];
      wr_data2 = wdata_i[2*WORD_WIDTH+:WORD_WIDTH];
      wr_data3 = wdata_i[3*WORD_WIDTH+:WORD_WIDTH];
    end
  end

  // RAM Bank 0 - Simple BRAM Template
  always_ff @(posedge clk_i) begin
    if (we0) begin
      ram0[wr_addr] <= wr_data0;
      rdata_q0 <= wr_data0;  // Write-first
    end else begin
      rdata_q0 <= ram0[word_addr];
    end
  end

  // RAM Bank 1 - Simple BRAM Template
  always_ff @(posedge clk_i) begin
    if (we1) begin
      ram1[wr_addr] <= wr_data1;
      rdata_q1 <= wr_data1;  // Write-first
    end else begin
      rdata_q1 <= ram1[word_addr];
    end
  end

  // RAM Bank 2 - Simple BRAM Template
  always_ff @(posedge clk_i) begin
    if (we2) begin
      ram2[wr_addr] <= wr_data2;
      rdata_q2 <= wr_data2;  // Write-first
    end else begin
      rdata_q2 <= ram2[word_addr];
    end
  end

  // RAM Bank 3 - Simple BRAM Template
  always_ff @(posedge clk_i) begin
    if (we3) begin
      ram3[wr_addr] <= wr_data3;
      rdata_q3 <= wr_data3;  // Write-first
    end else begin
      rdata_q3 <= ram3[word_addr];
    end
  end

  // Concatenate separate output registers
  assign rdata_o = {rdata_q3, rdata_q2, rdata_q1, rdata_q0};

  // ==========================================================================
  // Programming Module Instance
  // ==========================================================================
  ram_programmer #(
      .CLK_FREQ    (CPU_CLK),
      .BAUD_RATE   (PROG_BAUD_RATE),
      .MAGIC_SEQ   (PROGRAM_SEQUENCE),
      .SEQ_LENGTH  (PROGRAM_SEQUENCE_LEN),
      .BREAK_CYCLES(1_000_000)
  ) i_programmer (
      .clk_i         (clk_i),
      .rst_ni        (rst_ni),
      .uart_rx_i     (ram_prog_rx_i),
      .prog_addr_o   (prog_addr),
      .prog_data_o   (prog_data),
      .prog_valid_o  (prog_valid),
      .prog_mode_o   (prog_mode),
      .system_reset_o(prog_sys_rst)
  );

  // ==========================================================================
  // Output Assignments
  // ==========================================================================
  assign system_reset_o  = prog_sys_rst;
  assign prog_mode_led_o = prog_mode;

endmodule
