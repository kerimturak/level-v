/*
Copyright (c) 2025 Kerim TURAK

Permission is granted to use, copy, modify, and distribute this software for any purpose,
with or without fee, provided that the above notice appears in all copies.

THE SOFTWARE IS PROVIDED "AS IS" WITHOUT ANY WARRANTY OF ANY KIND.

================================================================================
VGA Character ROM (8x16 Font)
================================================================================
Description:
  8x16 pixel character ROM for VGA text mode.
  Contains ASCII characters 0-255.
  Each character is 16 bytes (16 rows of 8 pixels).

  Address = (char_code * 16) + row
  Data = 8-bit row bitmap (MSB = leftmost pixel)

  This is a subset containing printable ASCII (32-127).
  Extended characters can be added for code pages.
================================================================================
*/

`timescale 1ns / 1ps

module vga_char_rom (
    input  logic        clk_i,
    input  logic [11:0] addr_i,  // Character address (char * 16 + row)
    output logic [ 7:0] data_o
);

  // 256 characters * 16 rows = 4096 bytes
  logic [7:0] rom[4096];

  // Synchronous ROM read
  always_ff @(posedge clk_i) begin
    data_o <= rom[addr_i];
  end

  // Initialize ROM with 8x16 font
  initial begin
    // Clear all
    for (int i = 0; i < 4096; i++) begin
      rom[i] = 8'h00;
    end

    // Space (32)
    // All zeros - already initialized

    // ! (33)
    rom[33*16+1]   = 8'b00011000;
    rom[33*16+2]   = 8'b00111100;
    rom[33*16+3]   = 8'b00111100;
    rom[33*16+4]   = 8'b00111100;
    rom[33*16+5]   = 8'b00011000;
    rom[33*16+6]   = 8'b00011000;
    rom[33*16+7]   = 8'b00011000;
    rom[33*16+8]   = 8'b00000000;
    rom[33*16+9]   = 8'b00011000;
    rom[33*16+10]  = 8'b00011000;

    // " (34)
    rom[34*16+1]   = 8'b01100110;
    rom[34*16+2]   = 8'b01100110;
    rom[34*16+3]   = 8'b01100110;
    rom[34*16+4]   = 8'b00100100;

    // # (35)
    rom[35*16+2]   = 8'b01101100;
    rom[35*16+3]   = 8'b01101100;
    rom[35*16+4]   = 8'b11111110;
    rom[35*16+5]   = 8'b01101100;
    rom[35*16+6]   = 8'b11111110;
    rom[35*16+7]   = 8'b01101100;
    rom[35*16+8]   = 8'b01101100;

    // 0 (48)
    rom[48*16+2]   = 8'b01111100;
    rom[48*16+3]   = 8'b11000110;
    rom[48*16+4]   = 8'b11001110;
    rom[48*16+5]   = 8'b11011110;
    rom[48*16+6]   = 8'b11110110;
    rom[48*16+7]   = 8'b11100110;
    rom[48*16+8]   = 8'b11000110;
    rom[48*16+9]   = 8'b01111100;

    // 1 (49)
    rom[49*16+2]   = 8'b00011000;
    rom[49*16+3]   = 8'b00111000;
    rom[49*16+4]   = 8'b01111000;
    rom[49*16+5]   = 8'b00011000;
    rom[49*16+6]   = 8'b00011000;
    rom[49*16+7]   = 8'b00011000;
    rom[49*16+8]   = 8'b00011000;
    rom[49*16+9]   = 8'b01111110;

    // 2 (50)
    rom[50*16+2]   = 8'b01111100;
    rom[50*16+3]   = 8'b11000110;
    rom[50*16+4]   = 8'b00000110;
    rom[50*16+5]   = 8'b00001100;
    rom[50*16+6]   = 8'b00011000;
    rom[50*16+7]   = 8'b00110000;
    rom[50*16+8]   = 8'b01100000;
    rom[50*16+9]   = 8'b11111110;

    // 3 (51)
    rom[51*16+2]   = 8'b01111100;
    rom[51*16+3]   = 8'b11000110;
    rom[51*16+4]   = 8'b00000110;
    rom[51*16+5]   = 8'b00111100;
    rom[51*16+6]   = 8'b00000110;
    rom[51*16+7]   = 8'b00000110;
    rom[51*16+8]   = 8'b11000110;
    rom[51*16+9]   = 8'b01111100;

    // 4 (52)
    rom[52*16+2]   = 8'b00001100;
    rom[52*16+3]   = 8'b00011100;
    rom[52*16+4]   = 8'b00111100;
    rom[52*16+5]   = 8'b01101100;
    rom[52*16+6]   = 8'b11001100;
    rom[52*16+7]   = 8'b11111110;
    rom[52*16+8]   = 8'b00001100;
    rom[52*16+9]   = 8'b00011110;

    // 5 (53)
    rom[53*16+2]   = 8'b11111110;
    rom[53*16+3]   = 8'b11000000;
    rom[53*16+4]   = 8'b11000000;
    rom[53*16+5]   = 8'b11111100;
    rom[53*16+6]   = 8'b00000110;
    rom[53*16+7]   = 8'b00000110;
    rom[53*16+8]   = 8'b11000110;
    rom[53*16+9]   = 8'b01111100;

    // 6 (54)
    rom[54*16+2]   = 8'b00111100;
    rom[54*16+3]   = 8'b01100000;
    rom[54*16+4]   = 8'b11000000;
    rom[54*16+5]   = 8'b11111100;
    rom[54*16+6]   = 8'b11000110;
    rom[54*16+7]   = 8'b11000110;
    rom[54*16+8]   = 8'b11000110;
    rom[54*16+9]   = 8'b01111100;

    // 7 (55)
    rom[55*16+2]   = 8'b11111110;
    rom[55*16+3]   = 8'b11000110;
    rom[55*16+4]   = 8'b00000110;
    rom[55*16+5]   = 8'b00001100;
    rom[55*16+6]   = 8'b00011000;
    rom[55*16+7]   = 8'b00110000;
    rom[55*16+8]   = 8'b00110000;
    rom[55*16+9]   = 8'b00110000;

    // 8 (56)
    rom[56*16+2]   = 8'b01111100;
    rom[56*16+3]   = 8'b11000110;
    rom[56*16+4]   = 8'b11000110;
    rom[56*16+5]   = 8'b01111100;
    rom[56*16+6]   = 8'b11000110;
    rom[56*16+7]   = 8'b11000110;
    rom[56*16+8]   = 8'b11000110;
    rom[56*16+9]   = 8'b01111100;

    // 9 (57)
    rom[57*16+2]   = 8'b01111100;
    rom[57*16+3]   = 8'b11000110;
    rom[57*16+4]   = 8'b11000110;
    rom[57*16+5]   = 8'b01111110;
    rom[57*16+6]   = 8'b00000110;
    rom[57*16+7]   = 8'b00000110;
    rom[57*16+8]   = 8'b00001100;
    rom[57*16+9]   = 8'b01111000;

    // A (65)
    rom[65*16+2]   = 8'b00010000;
    rom[65*16+3]   = 8'b00111000;
    rom[65*16+4]   = 8'b01101100;
    rom[65*16+5]   = 8'b11000110;
    rom[65*16+6]   = 8'b11000110;
    rom[65*16+7]   = 8'b11111110;
    rom[65*16+8]   = 8'b11000110;
    rom[65*16+9]   = 8'b11000110;

    // B (66)
    rom[66*16+2]   = 8'b11111100;
    rom[66*16+3]   = 8'b01100110;
    rom[66*16+4]   = 8'b01100110;
    rom[66*16+5]   = 8'b01111100;
    rom[66*16+6]   = 8'b01100110;
    rom[66*16+7]   = 8'b01100110;
    rom[66*16+8]   = 8'b01100110;
    rom[66*16+9]   = 8'b11111100;

    // C (67)
    rom[67*16+2]   = 8'b00111100;
    rom[67*16+3]   = 8'b01100110;
    rom[67*16+4]   = 8'b11000000;
    rom[67*16+5]   = 8'b11000000;
    rom[67*16+6]   = 8'b11000000;
    rom[67*16+7]   = 8'b11000000;
    rom[67*16+8]   = 8'b01100110;
    rom[67*16+9]   = 8'b00111100;

    // D (68)
    rom[68*16+2]   = 8'b11111000;
    rom[68*16+3]   = 8'b01101100;
    rom[68*16+4]   = 8'b01100110;
    rom[68*16+5]   = 8'b01100110;
    rom[68*16+6]   = 8'b01100110;
    rom[68*16+7]   = 8'b01100110;
    rom[68*16+8]   = 8'b01101100;
    rom[68*16+9]   = 8'b11111000;

    // E (69)
    rom[69*16+2]   = 8'b11111110;
    rom[69*16+3]   = 8'b01100010;
    rom[69*16+4]   = 8'b01101000;
    rom[69*16+5]   = 8'b01111000;
    rom[69*16+6]   = 8'b01101000;
    rom[69*16+7]   = 8'b01100000;
    rom[69*16+8]   = 8'b01100010;
    rom[69*16+9]   = 8'b11111110;

    // F (70)
    rom[70*16+2]   = 8'b11111110;
    rom[70*16+3]   = 8'b01100010;
    rom[70*16+4]   = 8'b01101000;
    rom[70*16+5]   = 8'b01111000;
    rom[70*16+6]   = 8'b01101000;
    rom[70*16+7]   = 8'b01100000;
    rom[70*16+8]   = 8'b01100000;
    rom[70*16+9]   = 8'b11110000;

    // G (71)
    rom[71*16+2]   = 8'b00111100;
    rom[71*16+3]   = 8'b01100110;
    rom[71*16+4]   = 8'b11000000;
    rom[71*16+5]   = 8'b11000000;
    rom[71*16+6]   = 8'b11001110;
    rom[71*16+7]   = 8'b11000110;
    rom[71*16+8]   = 8'b01100110;
    rom[71*16+9]   = 8'b00111110;

    // H (72)
    rom[72*16+2]   = 8'b11000110;
    rom[72*16+3]   = 8'b11000110;
    rom[72*16+4]   = 8'b11000110;
    rom[72*16+5]   = 8'b11111110;
    rom[72*16+6]   = 8'b11000110;
    rom[72*16+7]   = 8'b11000110;
    rom[72*16+8]   = 8'b11000110;
    rom[72*16+9]   = 8'b11000110;

    // I (73)
    rom[73*16+2]   = 8'b00111100;
    rom[73*16+3]   = 8'b00011000;
    rom[73*16+4]   = 8'b00011000;
    rom[73*16+5]   = 8'b00011000;
    rom[73*16+6]   = 8'b00011000;
    rom[73*16+7]   = 8'b00011000;
    rom[73*16+8]   = 8'b00011000;
    rom[73*16+9]   = 8'b00111100;

    // J (74)
    rom[74*16+2]   = 8'b00011110;
    rom[74*16+3]   = 8'b00001100;
    rom[74*16+4]   = 8'b00001100;
    rom[74*16+5]   = 8'b00001100;
    rom[74*16+6]   = 8'b00001100;
    rom[74*16+7]   = 8'b11001100;
    rom[74*16+8]   = 8'b11001100;
    rom[74*16+9]   = 8'b01111000;

    // K (75)
    rom[75*16+2]   = 8'b11100110;
    rom[75*16+3]   = 8'b01100110;
    rom[75*16+4]   = 8'b01101100;
    rom[75*16+5]   = 8'b01111000;
    rom[75*16+6]   = 8'b01101100;
    rom[75*16+7]   = 8'b01100110;
    rom[75*16+8]   = 8'b01100110;
    rom[75*16+9]   = 8'b11100110;

    // L (76)
    rom[76*16+2]   = 8'b11110000;
    rom[76*16+3]   = 8'b01100000;
    rom[76*16+4]   = 8'b01100000;
    rom[76*16+5]   = 8'b01100000;
    rom[76*16+6]   = 8'b01100000;
    rom[76*16+7]   = 8'b01100000;
    rom[76*16+8]   = 8'b01100010;
    rom[76*16+9]   = 8'b11111110;

    // M (77)
    rom[77*16+2]   = 8'b11000110;
    rom[77*16+3]   = 8'b11101110;
    rom[77*16+4]   = 8'b11111110;
    rom[77*16+5]   = 8'b11111110;
    rom[77*16+6]   = 8'b11010110;
    rom[77*16+7]   = 8'b11000110;
    rom[77*16+8]   = 8'b11000110;
    rom[77*16+9]   = 8'b11000110;

    // N (78)
    rom[78*16+2]   = 8'b11000110;
    rom[78*16+3]   = 8'b11100110;
    rom[78*16+4]   = 8'b11110110;
    rom[78*16+5]   = 8'b11111110;
    rom[78*16+6]   = 8'b11011110;
    rom[78*16+7]   = 8'b11001110;
    rom[78*16+8]   = 8'b11000110;
    rom[78*16+9]   = 8'b11000110;

    // O (79)
    rom[79*16+2]   = 8'b01111100;
    rom[79*16+3]   = 8'b11000110;
    rom[79*16+4]   = 8'b11000110;
    rom[79*16+5]   = 8'b11000110;
    rom[79*16+6]   = 8'b11000110;
    rom[79*16+7]   = 8'b11000110;
    rom[79*16+8]   = 8'b11000110;
    rom[79*16+9]   = 8'b01111100;

    // P (80)
    rom[80*16+2]   = 8'b11111100;
    rom[80*16+3]   = 8'b01100110;
    rom[80*16+4]   = 8'b01100110;
    rom[80*16+5]   = 8'b01100110;
    rom[80*16+6]   = 8'b01111100;
    rom[80*16+7]   = 8'b01100000;
    rom[80*16+8]   = 8'b01100000;
    rom[80*16+9]   = 8'b11110000;

    // Q (81)
    rom[81*16+2]   = 8'b01111100;
    rom[81*16+3]   = 8'b11000110;
    rom[81*16+4]   = 8'b11000110;
    rom[81*16+5]   = 8'b11000110;
    rom[81*16+6]   = 8'b11000110;
    rom[81*16+7]   = 8'b11010110;
    rom[81*16+8]   = 8'b11011110;
    rom[81*16+9]   = 8'b01111100;
    rom[81*16+10]  = 8'b00001110;

    // R (82)
    rom[82*16+2]   = 8'b11111100;
    rom[82*16+3]   = 8'b01100110;
    rom[82*16+4]   = 8'b01100110;
    rom[82*16+5]   = 8'b01100110;
    rom[82*16+6]   = 8'b01111100;
    rom[82*16+7]   = 8'b01101100;
    rom[82*16+8]   = 8'b01100110;
    rom[82*16+9]   = 8'b11100110;

    // S (83)
    rom[83*16+2]   = 8'b01111100;
    rom[83*16+3]   = 8'b11000110;
    rom[83*16+4]   = 8'b01100000;
    rom[83*16+5]   = 8'b00111000;
    rom[83*16+6]   = 8'b00001100;
    rom[83*16+7]   = 8'b00000110;
    rom[83*16+8]   = 8'b11000110;
    rom[83*16+9]   = 8'b01111100;

    // T (84)
    rom[84*16+2]   = 8'b01111110;
    rom[84*16+3]   = 8'b01111110;
    rom[84*16+4]   = 8'b01011010;
    rom[84*16+5]   = 8'b00011000;
    rom[84*16+6]   = 8'b00011000;
    rom[84*16+7]   = 8'b00011000;
    rom[84*16+8]   = 8'b00011000;
    rom[84*16+9]   = 8'b00111100;

    // U (85)
    rom[85*16+2]   = 8'b11000110;
    rom[85*16+3]   = 8'b11000110;
    rom[85*16+4]   = 8'b11000110;
    rom[85*16+5]   = 8'b11000110;
    rom[85*16+6]   = 8'b11000110;
    rom[85*16+7]   = 8'b11000110;
    rom[85*16+8]   = 8'b11000110;
    rom[85*16+9]   = 8'b01111100;

    // V (86)
    rom[86*16+2]   = 8'b11000110;
    rom[86*16+3]   = 8'b11000110;
    rom[86*16+4]   = 8'b11000110;
    rom[86*16+5]   = 8'b11000110;
    rom[86*16+6]   = 8'b11000110;
    rom[86*16+7]   = 8'b01101100;
    rom[86*16+8]   = 8'b00111000;
    rom[86*16+9]   = 8'b00010000;

    // W (87)
    rom[87*16+2]   = 8'b11000110;
    rom[87*16+3]   = 8'b11000110;
    rom[87*16+4]   = 8'b11000110;
    rom[87*16+5]   = 8'b11010110;
    rom[87*16+6]   = 8'b11111110;
    rom[87*16+7]   = 8'b11111110;
    rom[87*16+8]   = 8'b11101110;
    rom[87*16+9]   = 8'b11000110;

    // X (88)
    rom[88*16+2]   = 8'b11000110;
    rom[88*16+3]   = 8'b11000110;
    rom[88*16+4]   = 8'b01101100;
    rom[88*16+5]   = 8'b00111000;
    rom[88*16+6]   = 8'b00111000;
    rom[88*16+7]   = 8'b01101100;
    rom[88*16+8]   = 8'b11000110;
    rom[88*16+9]   = 8'b11000110;

    // Y (89)
    rom[89*16+2]   = 8'b01100110;
    rom[89*16+3]   = 8'b01100110;
    rom[89*16+4]   = 8'b01100110;
    rom[89*16+5]   = 8'b00111100;
    rom[89*16+6]   = 8'b00011000;
    rom[89*16+7]   = 8'b00011000;
    rom[89*16+8]   = 8'b00011000;
    rom[89*16+9]   = 8'b00111100;

    // Z (90)
    rom[90*16+2]   = 8'b11111110;
    rom[90*16+3]   = 8'b11000110;
    rom[90*16+4]   = 8'b00001100;
    rom[90*16+5]   = 8'b00011000;
    rom[90*16+6]   = 8'b00110000;
    rom[90*16+7]   = 8'b01100000;
    rom[90*16+8]   = 8'b11000110;
    rom[90*16+9]   = 8'b11111110;

    // a (97)
    rom[97*16+4]   = 8'b01111000;
    rom[97*16+5]   = 8'b00001100;
    rom[97*16+6]   = 8'b01111100;
    rom[97*16+7]   = 8'b11001100;
    rom[97*16+8]   = 8'b11001100;
    rom[97*16+9]   = 8'b01110110;

    // b (98)
    rom[98*16+2]   = 8'b11100000;
    rom[98*16+3]   = 8'b01100000;
    rom[98*16+4]   = 8'b01100000;
    rom[98*16+5]   = 8'b01111100;
    rom[98*16+6]   = 8'b01100110;
    rom[98*16+7]   = 8'b01100110;
    rom[98*16+8]   = 8'b01100110;
    rom[98*16+9]   = 8'b11011100;

    // c (99)
    rom[99*16+4]   = 8'b01111100;
    rom[99*16+5]   = 8'b11000110;
    rom[99*16+6]   = 8'b11000000;
    rom[99*16+7]   = 8'b11000000;
    rom[99*16+8]   = 8'b11000110;
    rom[99*16+9]   = 8'b01111100;

    // d (100)
    rom[100*16+2]  = 8'b00011100;
    rom[100*16+3]  = 8'b00001100;
    rom[100*16+4]  = 8'b00001100;
    rom[100*16+5]  = 8'b01111100;
    rom[100*16+6]  = 8'b11001100;
    rom[100*16+7]  = 8'b11001100;
    rom[100*16+8]  = 8'b11001100;
    rom[100*16+9]  = 8'b01110110;

    // e (101)
    rom[101*16+4]  = 8'b01111100;
    rom[101*16+5]  = 8'b11000110;
    rom[101*16+6]  = 8'b11111110;
    rom[101*16+7]  = 8'b11000000;
    rom[101*16+8]  = 8'b11000110;
    rom[101*16+9]  = 8'b01111100;

    // f (102)
    rom[102*16+2]  = 8'b00111000;
    rom[102*16+3]  = 8'b01101100;
    rom[102*16+4]  = 8'b01100000;
    rom[102*16+5]  = 8'b11110000;
    rom[102*16+6]  = 8'b01100000;
    rom[102*16+7]  = 8'b01100000;
    rom[102*16+8]  = 8'b01100000;
    rom[102*16+9]  = 8'b11110000;

    // g (103)
    rom[103*16+4]  = 8'b01110110;
    rom[103*16+5]  = 8'b11001100;
    rom[103*16+6]  = 8'b11001100;
    rom[103*16+7]  = 8'b11001100;
    rom[103*16+8]  = 8'b01111100;
    rom[103*16+9]  = 8'b00001100;
    rom[103*16+10] = 8'b11001100;
    rom[103*16+11] = 8'b01111000;

    // h (104)
    rom[104*16+2]  = 8'b11100000;
    rom[104*16+3]  = 8'b01100000;
    rom[104*16+4]  = 8'b01100000;
    rom[104*16+5]  = 8'b01101100;
    rom[104*16+6]  = 8'b01110110;
    rom[104*16+7]  = 8'b01100110;
    rom[104*16+8]  = 8'b01100110;
    rom[104*16+9]  = 8'b11100110;

    // i (105)
    rom[105*16+2]  = 8'b00011000;
    rom[105*16+3]  = 8'b00000000;
    rom[105*16+4]  = 8'b00111000;
    rom[105*16+5]  = 8'b00011000;
    rom[105*16+6]  = 8'b00011000;
    rom[105*16+7]  = 8'b00011000;
    rom[105*16+8]  = 8'b00011000;
    rom[105*16+9]  = 8'b00111100;

    // j (106)
    rom[106*16+2]  = 8'b00000110;
    rom[106*16+3]  = 8'b00000000;
    rom[106*16+4]  = 8'b00001110;
    rom[106*16+5]  = 8'b00000110;
    rom[106*16+6]  = 8'b00000110;
    rom[106*16+7]  = 8'b00000110;
    rom[106*16+8]  = 8'b00000110;
    rom[106*16+9]  = 8'b01100110;
    rom[106*16+10] = 8'b01100110;
    rom[106*16+11] = 8'b00111100;

    // k (107)
    rom[107*16+2]  = 8'b11100000;
    rom[107*16+3]  = 8'b01100000;
    rom[107*16+4]  = 8'b01100110;
    rom[107*16+5]  = 8'b01101100;
    rom[107*16+6]  = 8'b01111000;
    rom[107*16+7]  = 8'b01101100;
    rom[107*16+8]  = 8'b01100110;
    rom[107*16+9]  = 8'b11100110;

    // l (108)
    rom[108*16+2]  = 8'b00111000;
    rom[108*16+3]  = 8'b00011000;
    rom[108*16+4]  = 8'b00011000;
    rom[108*16+5]  = 8'b00011000;
    rom[108*16+6]  = 8'b00011000;
    rom[108*16+7]  = 8'b00011000;
    rom[108*16+8]  = 8'b00011000;
    rom[108*16+9]  = 8'b00111100;

    // m (109)
    rom[109*16+4]  = 8'b11101100;
    rom[109*16+5]  = 8'b11111110;
    rom[109*16+6]  = 8'b11010110;
    rom[109*16+7]  = 8'b11010110;
    rom[109*16+8]  = 8'b11010110;
    rom[109*16+9]  = 8'b11000110;

    // n (110)
    rom[110*16+4]  = 8'b11011100;
    rom[110*16+5]  = 8'b01100110;
    rom[110*16+6]  = 8'b01100110;
    rom[110*16+7]  = 8'b01100110;
    rom[110*16+8]  = 8'b01100110;
    rom[110*16+9]  = 8'b01100110;

    // o (111)
    rom[111*16+4]  = 8'b01111100;
    rom[111*16+5]  = 8'b11000110;
    rom[111*16+6]  = 8'b11000110;
    rom[111*16+7]  = 8'b11000110;
    rom[111*16+8]  = 8'b11000110;
    rom[111*16+9]  = 8'b01111100;

    // p (112)
    rom[112*16+4]  = 8'b11011100;
    rom[112*16+5]  = 8'b01100110;
    rom[112*16+6]  = 8'b01100110;
    rom[112*16+7]  = 8'b01100110;
    rom[112*16+8]  = 8'b01111100;
    rom[112*16+9]  = 8'b01100000;
    rom[112*16+10] = 8'b01100000;
    rom[112*16+11] = 8'b11110000;

    // q (113)
    rom[113*16+4]  = 8'b01110110;
    rom[113*16+5]  = 8'b11001100;
    rom[113*16+6]  = 8'b11001100;
    rom[113*16+7]  = 8'b11001100;
    rom[113*16+8]  = 8'b01111100;
    rom[113*16+9]  = 8'b00001100;
    rom[113*16+10] = 8'b00001100;
    rom[113*16+11] = 8'b00011110;

    // r (114)
    rom[114*16+4]  = 8'b11011100;
    rom[114*16+5]  = 8'b01110110;
    rom[114*16+6]  = 8'b01100110;
    rom[114*16+7]  = 8'b01100000;
    rom[114*16+8]  = 8'b01100000;
    rom[114*16+9]  = 8'b11110000;

    // s (115)
    rom[115*16+4]  = 8'b01111100;
    rom[115*16+5]  = 8'b11000110;
    rom[115*16+6]  = 8'b01110000;
    rom[115*16+7]  = 8'b00011100;
    rom[115*16+8]  = 8'b11000110;
    rom[115*16+9]  = 8'b01111100;

    // t (116)
    rom[116*16+2]  = 8'b00010000;
    rom[116*16+3]  = 8'b00110000;
    rom[116*16+4]  = 8'b01111100;
    rom[116*16+5]  = 8'b00110000;
    rom[116*16+6]  = 8'b00110000;
    rom[116*16+7]  = 8'b00110000;
    rom[116*16+8]  = 8'b00110100;
    rom[116*16+9]  = 8'b00011000;

    // u (117)
    rom[117*16+4]  = 8'b11001100;
    rom[117*16+5]  = 8'b11001100;
    rom[117*16+6]  = 8'b11001100;
    rom[117*16+7]  = 8'b11001100;
    rom[117*16+8]  = 8'b11001100;
    rom[117*16+9]  = 8'b01110110;

    // v (118)
    rom[118*16+4]  = 8'b11001100;
    rom[118*16+5]  = 8'b11001100;
    rom[118*16+6]  = 8'b11001100;
    rom[118*16+7]  = 8'b11001100;
    rom[118*16+8]  = 8'b01111000;
    rom[118*16+9]  = 8'b00110000;

    // w (119)
    rom[119*16+4]  = 8'b11000110;
    rom[119*16+5]  = 8'b11000110;
    rom[119*16+6]  = 8'b11010110;
    rom[119*16+7]  = 8'b11111110;
    rom[119*16+8]  = 8'b11111110;
    rom[119*16+9]  = 8'b01101100;

    // x (120)
    rom[120*16+4]  = 8'b11000110;
    rom[120*16+5]  = 8'b01101100;
    rom[120*16+6]  = 8'b00111000;
    rom[120*16+7]  = 8'b00111000;
    rom[120*16+8]  = 8'b01101100;
    rom[120*16+9]  = 8'b11000110;

    // y (121)
    rom[121*16+4]  = 8'b11001100;
    rom[121*16+5]  = 8'b11001100;
    rom[121*16+6]  = 8'b11001100;
    rom[121*16+7]  = 8'b11001100;
    rom[121*16+8]  = 8'b01111100;
    rom[121*16+9]  = 8'b00001100;
    rom[121*16+10] = 8'b00011000;
    rom[121*16+11] = 8'b11110000;

    // z (122)
    rom[122*16+4]  = 8'b11111100;
    rom[122*16+5]  = 8'b10011000;
    rom[122*16+6]  = 8'b00110000;
    rom[122*16+7]  = 8'b01100000;
    rom[122*16+8]  = 8'b11000100;
    rom[122*16+9]  = 8'b11111100;
  end

endmodule
