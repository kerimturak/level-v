// ============================================================================
// Spike-like Commit Trace — Ceres RISC-V
// Engineer:  Kerim Turak
// ----------------------------------------------------------------------------
// Production order (Spike-compatible):
//   1. CSR write (wr_en_csr_i)
//   2. Memory write
//   3. Register writeback
//   4. No-write instruction
// 
// Enable with: +define+LOG_COMMIT
// ============================================================================

// Define SOC path based on top module name
`ifdef VERILATOR
  `define SOC $root.ceres_wrapper.i_soc
`else
  `define SOC tb_wrapper.ceres_wrapper.i_soc
`endif

`ifdef LOG_COMMIT

integer trace_fd;
string  trace_path;
string  test_name;
string  simulator;

// ============================================================================
// INITIAL (open trace file)
// ============================================================================
initial begin
  if (!$value$plusargs("simulator=%s", simulator))
    simulator = "default_simulator";

  if (!$value$plusargs("test_name=%s", test_name))
    test_name = "default_test";

  if (!$value$plusargs("trace_file=%s", trace_path))
    trace_path = $sformatf("/home/kerim/riscv_git/ceres-riscv/results/logs/%0s/%0s/commit_trace.log",
                            simulator, test_name);

  void'($system($sformatf("mkdir -p $(dirname %s)", trace_path)));

  trace_fd = $fopen(trace_path, "w");
  if (trace_fd == 0) begin
    $display("[ERROR] Failed to open trace file: %s", trace_path);
    $finish;
  end else begin
    $display("[COMMIT_LOG] Writing to: %s", trace_path);
  end
end

// ============================================================================
// MAIN TRACE LOGIC (Spike EXACT behavior)
// ============================================================================

always @(posedge clk_i) begin
  // Not: Reset sırasında dosyayı yeniden açmıyoruz - sadece initial'da açıldı
  if (rst_ni && !(stall_i inside {IMISS_STALL, DMISS_STALL, ALU_STALL, FENCEI_STALL} && !trap_active_i)) begin

    // Automatic variable for CSR WARL behavior:
    // - mstatus (0x300): MPP always 11 for M-mode only
    // - tselect (0x7A0): Read-only-zero (single trigger implementation)
    automatic logic [31:0] csr_log_value = (csr_idx_i == 12'h300) ? 
                                           (csr_wr_data_i | 32'h00001800) : 
                                           (csr_idx_i == 12'h7A0) ? 32'h0 :  // tselect: always 0
                                           csr_wr_data_i;

    // ============================================================
    // 1) SPIKE-STYLE: CSR + RD WRITE IN SAME INSTRUCTION (CSRRW / CSRRS / CSRRC)
    // ============================================================
    if ((instr_type_i inside {CSR_RW, CSR_RS, CSR_RC, CSR_RWI, CSR_RSI, CSR_RCI}) &&
        wr_en_csr_i && rf_rw_en_i && rd_addr_i != 0) begin

      // Format:
      // core 0: 3 PC (INST) x<rd> oldCSR  c<idx>_name newCSR
      $fwrite(trace_fd,
        "core   0: 3 0x%08h (0x%08h) x%0d 0x%08h c%0d_%s 0x%08h\n",
        pc_i,
        fe_tracer_i.inst,
        rd_addr_i,
        wb_data_o,                     // RD = OLD CSR
        csr_idx_i,
        csr_name(csr_idx_i),
        csr_log_value                  // CSR = NEW CSR with WARL applied
      );
    end

// ============================================================
// SPECIAL CASE — MRET implicit CSR writes
// Spike logs mstatus (0x300), mstatush (0x310), and tcontrol (0x7A5) on MRET.
// ============================================================
else if (instr_type_i == mret) begin : mret_commit

    // mstatus - apply WARL (MPP always 11)
    $fwrite(trace_fd,
      "core   0: 3 0x%08h (0x%08h) c%0d_mstatus 0x%08h ",
      pc_i, fe_tracer_i.inst,
      768,        // <<2 doğru
      csr_log_value
    );

    // mstatush
    $fwrite(trace_fd,
      "c%0d_mstatush 0x00000000 ",
      784         // <<2 doğru
    );

    // tcontrol - log actual value from CSR file
    $fwrite(trace_fd,
      "c%0d_tcontrol 0x%08h\n",
      1957,       // 0x7A5
      tcontrol_i
    );

    disable mret_commit;
end



    // ============================================================
    // 2) CSR WRITE ONLY (CSRWI, CSRRW x0,csr)
    // ============================================================
    else if (wr_en_csr_i) begin
      $fwrite(trace_fd,
        "core   0: 3 0x%08h (0x%08h) c%0d_%s 0x%08h\n",
        pc_i, fe_tracer_i.inst,
        csr_idx_i,
        csr_name(csr_idx_i),
        csr_log_value
      );
    end

    // ============================================================
    // 3) REGISTER WRITE ONLY (normal ALU, load result, jump-link, etc.)
    // ============================================================
    else if (instr_type_i inside {i_lb, i_lh, i_lw, i_lbu, i_lhu} && rd_addr_i != 0) begin
      automatic string spacing = (rd_addr_i < 10) ? "  " : " ";
      $fwrite(trace_fd,
        "core   0: 3 0x%08h (0x%08h) x%0d%s0x%08h mem 0x%08h\n",
        pc_i, fe_tracer_i.inst,
        rd_addr_i, spacing, wb_data_o,
        alu_result_i
      );
    end

    // Load to x0 - just log memory access without register write
    else if (instr_type_i inside {i_lb, i_lh, i_lw, i_lbu, i_lhu} && rd_addr_i == 0) begin
      $fwrite(trace_fd,
        "core   0: 3 0x%08h (0x%08h) mem 0x%08h\n",
        pc_i, fe_tracer_i.inst,
        alu_result_i
      );
    end

    else if (rf_rw_en_i && rd_addr_i != 0) begin
      automatic string spacing = (rd_addr_i < 10) ? "  " : " ";
      $fwrite(trace_fd,
        "core   0: 3 0x%08h (0x%08h) x%0d%s0x%08h\n",
        pc_i, fe_tracer_i.inst,
        rd_addr_i, spacing, wb_data_o
      );
    end

    // ============================================================
    // 4) MEMORY WRITE (store)
    // ============================================================
    else if (instr_type_i inside {s_sb, s_sh, s_sw}) begin
      automatic logic [31:0] wdata = write_data_i;

      case (rw_size_i)
        2'b01:
          $fwrite(trace_fd,
            "core   0: 3 0x%08h (0x%08h) mem 0x%08h 0x%02h\n",
            pc_i, fe_tracer_i.inst, alu_result_i, wdata[7:0]);

        2'b10:
          $fwrite(trace_fd,
            "core   0: 3 0x%08h (0x%08h) mem 0x%08h 0x%04h\n",
            pc_i, fe_tracer_i.inst, alu_result_i, wdata[15:0]);

        2'b11:
          $fwrite(trace_fd,
            "core   0: 3 0x%08h (0x%08h) mem 0x%08h 0x%08h\n",
            pc_i, fe_tracer_i.inst, alu_result_i, wdata[31:0]);
        default: ; // Do nothing for 2'b00
      endcase
    end

    // ============================================================
    // 5) NO-WRITE INSTRUCTION
    // ============================================================
    else begin
      $fwrite(trace_fd,
        "core   0: 3 0x%08h (0x%08h)\n",
        pc_i, fe_tracer_i.inst
      );
    end
  end
end

// Periyodik flush - her 65536 cycle'da bir buffer'ı diske yaz
// Reset-independent: initialization syntax kullanılıyor
logic [15:0] flush_counter = '0;
always @(posedge clk_i) begin
  if (rst_ni) begin
    flush_counter <= flush_counter + 1;
    if (flush_counter == 0 && trace_fd != 0) begin
      $fflush(trace_fd);
    end
  end
end

final begin
  if (trace_fd != 0) $fclose(trace_fd);
end

`endif // LOG_COMMIT

// ==========================================================
// PASS/FAIL Address Detector (from per-test addr.txt file)
// Disable with +no_addr plusarg
// This section is always active (not affected by FAST_SIM)
// ==========================================================

string addr_file;
`ifndef LOG_COMMIT
string test_name;  // Needed for legacy check below
`endif
logic [31:0] pass_addr, fail_addr;
logic addr_check_enabled;
integer addr_fd, r;

initial begin
  // Check if address checking is disabled
  if ($test$plusargs("no_addr")) begin
    $display("[INFO] Address checking disabled (+no_addr)");
    addr_check_enabled = 0;
    pass_addr = 32'h0;
    fail_addr = 32'h0;
  end
  // Dosya ismini +arg ile al: +addr_file=/path/to/test_addr.txt
  else if (!$value$plusargs("addr_file=%s", addr_file)) begin
    $display("[INFO] No +addr_file given. Skipping PASS/FAIL auto-stop.");
`ifdef NO_COMMIT_TRACE
    if (!$value$plusargs("test_name=%s", test_name)) test_name = "";
`endif
    if (test_name == "rv32ui-p-simple") begin
      pass_addr = 32'h8000013c;
      fail_addr = 32'h80000140;
      addr_check_enabled = 1;
    end else begin
      pass_addr = 32'h0;
      fail_addr = 32'h0;
      addr_check_enabled = 0;
    end
  end else begin
    addr_fd = $fopen(addr_file, "r");
    if (addr_fd == 0) begin
      $display("ERROR: cannot open %s", addr_file);
      pass_addr = 32'h0;
      fail_addr = 32'h0;
      addr_check_enabled = 0;
    end else begin
      r = $fscanf(addr_fd, "%h %h", pass_addr, fail_addr);
      $fclose(addr_fd);
      $display("Loaded PASS/FAIL addresses: PASS=0x%08h FAIL=0x%08h", pass_addr, fail_addr);
      addr_check_enabled = 1;
    end
  end
end

// Writeback veya memory stage içinde:
always_comb begin
  if (addr_check_enabled && pc_i == pass_addr && pass_addr != 32'h0) begin
    $display("🎯 PASS address reached at PC=0x%08h", pc_i);
    $finish;
  end else if (addr_check_enabled && pc_i == fail_addr && fail_addr != 32'h0) begin
    $display("FAIL address reached at PC=0x%08h", pc_i);
    $finish;
  end
end

task automatic check_pass_fail();
  if (addr_check_enabled && pass_addr != 32'h0 && pc_i == pass_addr) begin
    $display("PASS reached at PC=0x%08h", pc_i);
    $finish;
  end
  if (addr_check_enabled && fail_addr != 32'h0 && pc_i == fail_addr) begin
    $display("FAIL reached at PC=0x%08h", pc_i);
    $finish;
  end
endtask

// TOHOST check - only for riscv-tests (isa tests), not arch tests
// When addr_check_enabled is true, pass/fail is determined by PC addresses
// When addr_check_enabled is false, use TOHOST memory-mapped register
always @(posedge clk_i) begin
  automatic logic        we = wr_en_i;
  automatic logic        valid = `SOC.pipe4.dcache_valid;
  automatic logic [31:0] addr = `SOC.pipe4.alu_result;
  automatic logic [31:0] data = `SOC.pipe4.write_data;

  if (!addr_check_enabled && valid && we && addr == 32'h80001000) begin
    if (data == 32'h1) begin
      $display("🎉 TOHOST PASS");
      $finish;
    end else begin
      $display("❌ TOHOST FAIL (0x%08h)", data);
      $finish;
    end
  end
end
